module DLY3X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX5M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X8M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX12M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND4BBX1M (
	Y, 
	D, 
	C, 
	BN, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input BN;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X2M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA22X2M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFQX2M (
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFQX1M (
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4BBX1M (
	Y, 
	D, 
	C, 
	BN, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input BN;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI33X2M (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX1M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Mon Aug 26 23:41:23 2024
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN3_scan_rst;
   wire FE_PHN0_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC3_scan_rst (
	.Y(FE_PHN3_scan_rst),
	.A(FE_PHN0_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_scan_rst (
	.Y(FE_PHN0_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN3_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN5_scan_rst;
   wire FE_PHN2_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC5_scan_rst (
	.Y(FE_PHN5_scan_rst),
	.A(FE_PHN2_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_scan_rst (
	.Y(FE_PHN2_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X8M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN5_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN4_scan_rst;
   wire FE_PHN1_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC4_scan_rst (
	.Y(FE_PHN4_scan_rst),
	.A(FE_PHN1_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC1_scan_rst (
	.Y(FE_PHN1_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X8M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN4_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DATA_SYNC_BUS_WIDTH8_test_1 (
	CLK, 
	RST, 
	BUS_EN, 
	UN_SYNC_BUS, 
	EN_PULSE, 
	SYNC_BUS, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN8_SE, 
	FE_OFN9_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input BUS_EN;
   input [7:0] UN_SYNC_BUS;
   output EN_PULSE;
   output [7:0] SYNC_BUS;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN8_SE;
   input FE_OFN9_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire SYNC_BUS_EN;
   wire PULSE_GEN_OUT;
   wire N1;
   wire n3;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n23;
   wire [1:0] stages;

   assign test_so = stages[1] ;

   // Module instantiations
   SDFFRQX2M PULSE_GEN_OUT_reg (
	.SI(EN_PULSE),
	.SE(test_se),
	.RN(RST),
	.Q(PULSE_GEN_OUT),
	.D(SYNC_BUS_EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[7]  (
	.SI(SYNC_BUS[6]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(SYNC_BUS[7]),
	.D(n17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[6]  (
	.SI(SYNC_BUS[5]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(SYNC_BUS[6]),
	.D(n15),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[4]  (
	.SI(SYNC_BUS[3]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(SYNC_BUS[4]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M SYNC_BUS_EN_reg (
	.SI(PULSE_GEN_OUT),
	.SE(FE_OFN9_SE),
	.RN(RST),
	.Q(SYNC_BUS_EN),
	.D(stages[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[5]  (
	.SI(SYNC_BUS[4]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(SYNC_BUS[5]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[3]  (
	.SI(SYNC_BUS[2]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[3]),
	.D(n9),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[1]  (
	.SI(SYNC_BUS[0]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[1]),
	.D(n5),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[0]  (
	.SI(n23),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[0]),
	.D(n3),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_BUS_reg[2]  (
	.SI(SYNC_BUS[1]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_BUS[2]),
	.D(n7),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M EN_PULSE_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(EN_PULSE),
	.D(N1),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \stages_reg[0]  (
	.SI(SYNC_BUS[7]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(stages[0]),
	.D(BUS_EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \stages_reg[1]  (
	.SI(stages[0]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(stages[1]),
	.D(stages[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n23),
	.A(SYNC_BUS_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(N1),
	.B(n23),
	.A(PULSE_GEN_OUT), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n3),
	.B1(n23),
	.B0(SYNC_BUS[0]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n5),
	.B1(n23),
	.B0(SYNC_BUS[1]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n7),
	.B1(n23),
	.B0(SYNC_BUS[2]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n9),
	.B1(n23),
	.B0(SYNC_BUS[3]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n11),
	.B1(n23),
	.B0(SYNC_BUS[4]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n13),
	.B1(n23),
	.B0(SYNC_BUS[5]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n15),
	.B1(n23),
	.B0(SYNC_BUS[6]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n17),
	.B1(n23),
	.B0(SYNC_BUS[7]),
	.A1(SYNC_BUS_EN),
	.A0(UN_SYNC_BUS[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_CTRL_DATA_WIDTH8_ADDRESS_WIDTH4_FUN_WIDTH4_ALU_OUT_WIDTH16_test_1 (
	CLK, 
	RST, 
	RX_P_DATA, 
	RX_DATA_VALID, 
	RD_DATA, 
	RD_DATA_VALID, 
	ALU_OUT, 
	ALU_OUT_VALID, 
	FIFO_FULL, 
	ALU_FUN, 
	ALU_EN, 
	CLK_GATE_EN, 
	ADDRESS, 
	WR_EN, 
	RD_EN, 
	WR_DATA, 
	TX_P_Data, 
	TX_DATA_VALID, 
	CLK_DIV_EN, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN1_SYNC_REF_SCAN_RST, 
	FE_OFN7_SE, 
	FE_OFN8_SE, 
	REF_SCAN_CLK__L2_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] RX_P_DATA;
   input RX_DATA_VALID;
   input [7:0] RD_DATA;
   input RD_DATA_VALID;
   input [15:0] ALU_OUT;
   input ALU_OUT_VALID;
   input FIFO_FULL;
   output [3:0] ALU_FUN;
   output ALU_EN;
   output CLK_GATE_EN;
   output [3:0] ADDRESS;
   output WR_EN;
   output RD_EN;
   output [7:0] WR_DATA;
   output [7:0] TX_P_Data;
   output TX_DATA_VALID;
   output CLK_DIV_EN;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN1_SYNC_REF_SCAN_RST;
   input FE_OFN7_SE;
   input FE_OFN8_SE;
   input REF_SCAN_CLK__L2_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire FE_OFN5_ADDRESS_3_;
   wire FE_OFN4_ADDRESS_2_;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n29;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire [3:0] current_state;
   wire [3:0] next_state;

   assign test_so = n71 ;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC5_ADDRESS_3_ (
	.Y(ADDRESS[3]),
	.A(FE_OFN5_ADDRESS_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC4_ADDRESS_2_ (
	.Y(ADDRESS[2]),
	.A(FE_OFN4_ADDRESS_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[7]  (
	.SI(n153),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n48),
	.Q(n152),
	.D(n125),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[6]  (
	.SI(n154),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n49),
	.Q(n153),
	.D(n124),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[5]  (
	.SI(n155),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n50),
	.Q(n154),
	.D(n123),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[4]  (
	.SI(n156),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n51),
	.Q(n155),
	.D(n122),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[3]  (
	.SI(n157),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n52),
	.Q(n156),
	.D(n121),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[2]  (
	.SI(n158),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n53),
	.Q(n157),
	.D(n120),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[1]  (
	.SI(n159),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n54),
	.Q(n158),
	.D(n119),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[0]  (
	.SI(n160),
	.SE(test_se),
	.RN(RST),
	.QN(n55),
	.Q(n159),
	.D(n118),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[14]  (
	.SI(n146),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n41),
	.Q(n145),
	.D(n132),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[13]  (
	.SI(n147),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n42),
	.Q(n146),
	.D(n131),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[12]  (
	.SI(n148),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n43),
	.Q(n147),
	.D(n130),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[11]  (
	.SI(n149),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n44),
	.Q(n148),
	.D(n129),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[10]  (
	.SI(n150),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n45),
	.Q(n149),
	.D(n128),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[9]  (
	.SI(n151),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n46),
	.Q(n150),
	.D(n127),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[8]  (
	.SI(n152),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n47),
	.Q(n151),
	.D(n126),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ADDRESS_REG_reg[2]  (
	.SI(n162),
	.SE(test_se),
	.RN(RST),
	.QN(n37),
	.Q(n161),
	.D(n136),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ADDRESS_REG_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.QN(n39),
	.Q(n163),
	.D(n134),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ADDRESS_REG_reg[3]  (
	.SI(n161),
	.SE(test_se),
	.RN(RST),
	.QN(n36),
	.Q(n160),
	.D(n137),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ADDRESS_REG_reg[1]  (
	.SI(n163),
	.SE(test_se),
	.RN(RST),
	.QN(n38),
	.Q(n162),
	.D(n135),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n65),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[3]  (
	.SI(n69),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(current_state[3]),
	.D(next_state[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n70),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(n144),
	.SE(test_se),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \ALU_OUT_REG_reg[15]  (
	.SI(n145),
	.SE(FE_OFN8_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.QN(n40),
	.Q(n144),
	.D(n133),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U30 (
	.Y(FE_OFN4_ADDRESS_2_),
	.B1(n117),
	.B0(n37),
	.A1(n107),
	.A0(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U31 (
	.Y(n114),
	.D(current_state[2]),
	.C(current_state[0]),
	.B(n71),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n63),
	.A(WR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(WR_EN),
	.B(n106),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U34 (
	.Y(n117),
	.B(n72),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U35 (
	.Y(n111),
	.B(n32),
	.A(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n68),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n62),
	.A(n105), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n29),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n32),
	.A(FIFO_FULL), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U41 (
	.Y(n106),
	.C(n80),
	.B(n76),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n72),
	.A(RX_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U43 (
	.Y(n80),
	.C(n116),
	.B(n69),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U44 (
	.Y(WR_DATA[0]),
	.B(n109),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U45 (
	.Y(WR_DATA[1]),
	.B(n108),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U46 (
	.Y(WR_DATA[2]),
	.B(n107),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U47 (
	.Y(WR_DATA[3]),
	.B(n103),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(WR_DATA[5]),
	.B(n63),
	.A(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U49 (
	.Y(TX_DATA_VALID),
	.B0(n113),
	.A1(n115),
	.A0(FIFO_FULL), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U50 (
	.Y(n74),
	.B(n84),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U51 (
	.Y(n83),
	.B(n65),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U52 (
	.Y(RD_EN),
	.B(n72),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U53 (
	.Y(n115),
	.B(n114),
	.A(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U54 (
	.Y(n112),
	.B(n32),
	.A(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U55 (
	.Y(WR_DATA[4]),
	.B(n63),
	.A(n139), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U56 (
	.Y(WR_DATA[7]),
	.B(n63),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U57 (
	.Y(n99),
	.B(n71),
	.AN(n84), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U58 (
	.Y(n84),
	.B(n69),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U59 (
	.Y(n94),
	.B(RX_DATA_VALID),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U60 (
	.Y(next_state[1]),
	.C0(n81),
	.B0(n66),
	.A1(n80),
	.A0(RX_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U61 (
	.Y(n81),
	.C0(n83),
	.B0(n64),
	.A1(n82),
	.A0(RX_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U62 (
	.Y(n66),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U63 (
	.Y(n82),
	.B0(n76),
	.A1(n65),
	.A0(n84), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U64 (
	.Y(n105),
	.C(n99),
	.B(n65),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U65 (
	.Y(n102),
	.D(n103),
	.C(n138),
	.B(n142),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U66 (
	.Y(n97),
	.D(n138),
	.C(n142),
	.B(n139),
	.A(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U67 (
	.Y(n89),
	.B0(n76),
	.A1(n99),
	.A0(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U68 (
	.Y(n64),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U69 (
	.Y(next_state[3]),
	.B(n74),
	.A(ALU_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U70 (
	.Y(ALU_EN),
	.B(n95),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U71 (
	.Y(ALU_FUN[2]),
	.B(n107),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U72 (
	.Y(ALU_FUN[3]),
	.B(n103),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U73 (
	.Y(ALU_FUN[0]),
	.B(n109),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U74 (
	.Y(ALU_FUN[1]),
	.B(n108),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U76 (
	.Y(CLK_GATE_EN),
	.C(n115),
	.B(n68),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U77 (
	.Y(FE_OFN5_ADDRESS_3_),
	.B1(n117),
	.B0(n36),
	.A1(n103),
	.A0(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U78 (
	.Y(n110),
	.C(n69),
	.B(current_state[3]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U79 (
	.Y(n116),
	.B(current_state[3]),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U80 (
	.Y(n90),
	.C(current_state[0]),
	.B(n69),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U81 (
	.Y(n65),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U82 (
	.Y(n76),
	.B(current_state[0]),
	.A(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U83 (
	.Y(n69),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U84 (
	.Y(n98),
	.C(current_state[2]),
	.B(n65),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U86 (
	.Y(n70),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U87 (
	.Y(ADDRESS[0]),
	.C1(n109),
	.C0(n90),
	.B1(n117),
	.B0(n39),
	.A1(n98),
	.A0(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U88 (
	.Y(n79),
	.B1(n95),
	.B0(RX_DATA_VALID),
	.A2(n94),
	.A1(n93),
	.A0(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U89 (
	.Y(n92),
	.B(RX_P_DATA[0]),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U90 (
	.Y(n95),
	.C(current_state[2]),
	.B(n116),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U91 (
	.Y(n85),
	.C0(n67),
	.B0(n91),
	.A1(n90),
	.A0(RX_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U92 (
	.Y(n91),
	.D(n97),
	.C(n96),
	.B(RX_P_DATA[7]),
	.AN(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U93 (
	.Y(n67),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U94 (
	.Y(n96),
	.C(RX_P_DATA[2]),
	.B(RX_P_DATA[6]),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U95 (
	.Y(next_state[2]),
	.D(n77),
	.C(n76),
	.B(n75),
	.AN(RD_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U96 (
	.Y(n77),
	.C0(n64),
	.B0(n79),
	.A1(n33),
	.A0(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n33),
	.A(RD_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U98 (
	.Y(WR_DATA[6]),
	.B(n63),
	.AN(RX_P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U99 (
	.Y(TX_P_Data[0]),
	.C1(n61),
	.C0(n113),
	.B1(n112),
	.B0(n47),
	.A1(n111),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U100 (
	.Y(n61),
	.A(RD_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U101 (
	.Y(TX_P_Data[1]),
	.C1(n60),
	.C0(n113),
	.B1(n112),
	.B0(n46),
	.A1(n111),
	.A0(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U102 (
	.Y(n60),
	.A(RD_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U103 (
	.Y(TX_P_Data[2]),
	.C1(n59),
	.C0(n113),
	.B1(n112),
	.B0(n45),
	.A1(n111),
	.A0(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U104 (
	.Y(n59),
	.A(RD_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U105 (
	.Y(TX_P_Data[3]),
	.C1(n58),
	.C0(n113),
	.B1(n112),
	.B0(n44),
	.A1(n111),
	.A0(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n58),
	.A(RD_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U107 (
	.Y(TX_P_Data[4]),
	.C1(n57),
	.C0(n113),
	.B1(n112),
	.B0(n43),
	.A1(n111),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n57),
	.A(RD_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U109 (
	.Y(TX_P_Data[5]),
	.C1(n56),
	.C0(n113),
	.B1(n112),
	.B0(n42),
	.A1(n111),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U110 (
	.Y(n56),
	.A(RD_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U111 (
	.Y(TX_P_Data[6]),
	.C1(n35),
	.C0(n113),
	.B1(n112),
	.B0(n41),
	.A1(n111),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U112 (
	.Y(n35),
	.A(RD_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U113 (
	.Y(TX_P_Data[7]),
	.C1(n34),
	.C0(n113),
	.B1(n112),
	.B0(n40),
	.A1(n111),
	.A0(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U114 (
	.Y(n34),
	.A(RD_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U115 (
	.Y(n100),
	.B(current_state[0]),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U116 (
	.Y(n103),
	.B(RX_DATA_VALID),
	.A(RX_P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U117 (
	.Y(n113),
	.C(RD_DATA_VALID),
	.B(n32),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U118 (
	.Y(n78),
	.B(current_state[0]),
	.AN(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U119 (
	.Y(n107),
	.B(RX_DATA_VALID),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U120 (
	.Y(n108),
	.B(RX_DATA_VALID),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U121 (
	.Y(n109),
	.B(RX_DATA_VALID),
	.A(RX_P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U122 (
	.Y(n93),
	.D(n104),
	.C(RX_P_DATA[7]),
	.B(RX_P_DATA[3]),
	.A(RX_P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U123 (
	.Y(n104),
	.C(RX_P_DATA[1]),
	.B(RX_P_DATA[5]),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U124 (
	.Y(n71),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U125 (
	.Y(next_state[0]),
	.D(n88),
	.C(n87),
	.B(n86),
	.A(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U126 (
	.Y(n87),
	.D(n102),
	.C(n101),
	.B(n143),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U127 (
	.Y(n88),
	.C0(n85),
	.B1(RX_DATA_VALID),
	.B0(n64),
	.A1(n72),
	.A0(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U128 (
	.Y(n101),
	.C(RX_P_DATA[4]),
	.B(RX_P_DATA[6]),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U129 (
	.Y(n141),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U130 (
	.Y(ADDRESS[1]),
	.B1(n117),
	.B0(n38),
	.A1(n108),
	.A0(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U131 (
	.Y(n134),
	.B1(n39),
	.B0(n105),
	.A1(n62),
	.A0(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U132 (
	.Y(n135),
	.B1(n38),
	.B0(n105),
	.A1(n62),
	.A0(n142), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U133 (
	.Y(n136),
	.B1(n37),
	.B0(n105),
	.A1(n62),
	.A0(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U134 (
	.Y(n137),
	.B1(n36),
	.B0(n105),
	.A1(n62),
	.A0(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U135 (
	.Y(n86),
	.C(ALU_OUT_VALID),
	.B(n65),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n118),
	.B1(n55),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n119),
	.B1(n54),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n120),
	.B1(n53),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n121),
	.B1(n52),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n122),
	.B1(n51),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n123),
	.B1(n50),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n124),
	.B1(n49),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n125),
	.B1(n48),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n126),
	.B1(n47),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n127),
	.B1(n46),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n128),
	.B1(n45),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n129),
	.B1(n44),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n130),
	.B1(n43),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U149 (
	.Y(n131),
	.B1(n42),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U150 (
	.Y(n132),
	.B1(n41),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U151 (
	.Y(n133),
	.B1(n40),
	.B0(n29),
	.A1N(n29),
	.A0N(ALU_OUT[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U152 (
	.Y(n142),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U153 (
	.Y(n138),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U154 (
	.Y(n143),
	.A(RX_P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U155 (
	.Y(n139),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U156 (
	.Y(n73),
	.A(RX_P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U157 (
	.Y(n75),
	.D(RX_P_DATA[4]),
	.C(RX_P_DATA[0]),
	.B(n94),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U158 (
	.Y(n140),
	.A(RX_P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(CLK_DIV_EN),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_NUM_STAGES2_test_0 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [1:0] stages;

   assign test_so = stages[1] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M SYNC_RST_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(stages[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \stages_reg[0]  (
	.SI(SYNC_RST),
	.SE(test_se),
	.RN(RST),
	.Q(stages[0]),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \stages_reg[1]  (
	.SI(stages[0]),
	.SE(test_se),
	.RN(RST),
	.Q(stages[1]),
	.D(stages[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_NUM_STAGES2_test_1 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [1:0] stages;

   assign test_so = stages[1] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M SYNC_RST_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(stages[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \stages_reg[0]  (
	.SI(SYNC_RST),
	.SE(test_se),
	.RN(RST),
	.Q(stages[0]),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \stages_reg[1]  (
	.SI(stages[0]),
	.SE(test_se),
	.RN(RST),
	.Q(stages[1]),
	.D(stages[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Reg_File_DATA_WIDTH8_DEPTH16_ADDRESS_WIDTH4_test_1 (
	CLK, 
	RST, 
	WR_DATA, 
	ADDRESS, 
	WR_EN, 
	RD_EN, 
	RD_DATA, 
	RD_DATA_VALID, 
	REG_0, 
	REG_1, 
	REG_2, 
	REG_3, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN0_SYNC_REF_SCAN_RST, 
	FE_OFN1_SYNC_REF_SCAN_RST, 
	FE_OFN7_SE, 
	REF_SCAN_CLK__L2_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] WR_DATA;
   input [3:0] ADDRESS;
   input WR_EN;
   input RD_EN;
   output [7:0] RD_DATA;
   output RD_DATA_VALID;
   output [7:0] REG_0;
   output [7:0] REG_1;
   output [7:0] REG_2;
   output [7:0] REG_3;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN0_SYNC_REF_SCAN_RST;
   input FE_OFN1_SYNC_REF_SCAN_RST;
   input FE_OFN7_SE;
   input REF_SCAN_CLK__L2_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN13_SE;
   wire FE_OFN11_SE;
   wire FE_OFN2_SYNC_REF_SCAN_RST;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire \REG[15][7] ;
   wire \REG[15][6] ;
   wire \REG[15][5] ;
   wire \REG[15][4] ;
   wire \REG[15][3] ;
   wire \REG[15][2] ;
   wire \REG[15][1] ;
   wire \REG[15][0] ;
   wire \REG[14][7] ;
   wire \REG[14][6] ;
   wire \REG[14][5] ;
   wire \REG[14][4] ;
   wire \REG[14][3] ;
   wire \REG[14][2] ;
   wire \REG[14][1] ;
   wire \REG[14][0] ;
   wire \REG[13][7] ;
   wire \REG[13][6] ;
   wire \REG[13][5] ;
   wire \REG[13][4] ;
   wire \REG[13][3] ;
   wire \REG[13][2] ;
   wire \REG[13][1] ;
   wire \REG[13][0] ;
   wire \REG[12][7] ;
   wire \REG[12][6] ;
   wire \REG[12][5] ;
   wire \REG[12][4] ;
   wire \REG[12][3] ;
   wire \REG[12][2] ;
   wire \REG[12][1] ;
   wire \REG[12][0] ;
   wire \REG[11][7] ;
   wire \REG[11][6] ;
   wire \REG[11][5] ;
   wire \REG[11][4] ;
   wire \REG[11][3] ;
   wire \REG[11][2] ;
   wire \REG[11][1] ;
   wire \REG[11][0] ;
   wire \REG[10][7] ;
   wire \REG[10][6] ;
   wire \REG[10][5] ;
   wire \REG[10][4] ;
   wire \REG[10][3] ;
   wire \REG[10][2] ;
   wire \REG[10][1] ;
   wire \REG[10][0] ;
   wire \REG[9][7] ;
   wire \REG[9][6] ;
   wire \REG[9][5] ;
   wire \REG[9][4] ;
   wire \REG[9][3] ;
   wire \REG[9][2] ;
   wire \REG[9][1] ;
   wire \REG[9][0] ;
   wire \REG[8][7] ;
   wire \REG[8][6] ;
   wire \REG[8][5] ;
   wire \REG[8][4] ;
   wire \REG[8][3] ;
   wire \REG[8][2] ;
   wire \REG[8][1] ;
   wire \REG[8][0] ;
   wire \REG[7][7] ;
   wire \REG[7][6] ;
   wire \REG[7][5] ;
   wire \REG[7][4] ;
   wire \REG[7][3] ;
   wire \REG[7][2] ;
   wire \REG[7][1] ;
   wire \REG[7][0] ;
   wire \REG[6][7] ;
   wire \REG[6][6] ;
   wire \REG[6][5] ;
   wire \REG[6][4] ;
   wire \REG[6][3] ;
   wire \REG[6][2] ;
   wire \REG[6][1] ;
   wire \REG[6][0] ;
   wire \REG[5][7] ;
   wire \REG[5][6] ;
   wire \REG[5][5] ;
   wire \REG[5][4] ;
   wire \REG[5][3] ;
   wire \REG[5][2] ;
   wire \REG[5][1] ;
   wire \REG[5][0] ;
   wire \REG[4][7] ;
   wire \REG[4][6] ;
   wire \REG[4][5] ;
   wire \REG[4][4] ;
   wire \REG[4][3] ;
   wire \REG[4][2] ;
   wire \REG[4][1] ;
   wire \REG[4][0] ;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n336;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;

   assign N11 = ADDRESS[0] ;
   assign N12 = ADDRESS[1] ;
   assign N13 = ADDRESS[2] ;
   assign N14 = ADDRESS[3] ;
   assign test_so2 = \REG[15][7]  ;
   assign test_so1 = \REG[14][1]  ;

   // Module instantiations
   BUFX4M FE_OFC13_SE (
	.Y(FE_OFN13_SE),
	.A(FE_OFN11_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC11_SE (
	.Y(FE_OFN11_SE),
	.A(FE_OFN7_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC2_SYNC_REF_SCAN_RST (
	.Y(FE_OFN2_SYNC_REF_SCAN_RST),
	.A(FE_OFN0_SYNC_REF_SCAN_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][7]  (
	.SI(\REG[13][6] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][7] ),
	.D(n297),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][6]  (
	.SI(\REG[13][5] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][6] ),
	.D(n296),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][5]  (
	.SI(\REG[13][4] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][5] ),
	.D(n295),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][4]  (
	.SI(\REG[13][3] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][4] ),
	.D(n294),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][3]  (
	.SI(\REG[13][2] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][3] ),
	.D(n293),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][2]  (
	.SI(\REG[13][1] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][2] ),
	.D(n292),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][1]  (
	.SI(\REG[13][0] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][1] ),
	.D(n291),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[13][0]  (
	.SI(\REG[12][7] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[13][0] ),
	.D(n290),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][7]  (
	.SI(\REG[9][6] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[9][7] ),
	.D(n265),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][6]  (
	.SI(\REG[9][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[9][6] ),
	.D(n264),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][5]  (
	.SI(\REG[9][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[9][5] ),
	.D(n263),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][4]  (
	.SI(\REG[9][3] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[9][4] ),
	.D(n262),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][3]  (
	.SI(\REG[9][2] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[9][3] ),
	.D(n261),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][2]  (
	.SI(\REG[9][1] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[9][2] ),
	.D(n260),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][1]  (
	.SI(\REG[9][0] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[9][1] ),
	.D(n259),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[9][0]  (
	.SI(\REG[8][7] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[9][0] ),
	.D(n258),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][7]  (
	.SI(\REG[5][6] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[5][7] ),
	.D(n233),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][6]  (
	.SI(\REG[5][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[5][6] ),
	.D(n232),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][5]  (
	.SI(\REG[5][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[5][5] ),
	.D(n231),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][4]  (
	.SI(\REG[5][3] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[5][4] ),
	.D(n230),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][3]  (
	.SI(\REG[5][2] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[5][3] ),
	.D(n229),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][2]  (
	.SI(\REG[5][1] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[5][2] ),
	.D(n228),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][1]  (
	.SI(\REG[5][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[5][1] ),
	.D(n227),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5][0]  (
	.SI(\REG[4][7] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[5][0] ),
	.D(n226),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][7]  (
	.SI(\REG[15][6] ),
	.SE(test_se),
	.RN(RST),
	.Q(\REG[15][7] ),
	.D(n313),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][6]  (
	.SI(\REG[15][5] ),
	.SE(test_se),
	.RN(RST),
	.Q(\REG[15][6] ),
	.D(n312),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][5]  (
	.SI(\REG[15][4] ),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(\REG[15][5] ),
	.D(n311),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][4]  (
	.SI(\REG[15][3] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[15][4] ),
	.D(n310),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][3]  (
	.SI(\REG[15][2] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[15][3] ),
	.D(n309),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][2]  (
	.SI(\REG[15][1] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[15][2] ),
	.D(n308),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][1]  (
	.SI(\REG[15][0] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[15][1] ),
	.D(n307),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[15][0]  (
	.SI(\REG[14][7] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[15][0] ),
	.D(n306),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][7]  (
	.SI(\REG[11][6] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[11][7] ),
	.D(n281),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][6]  (
	.SI(\REG[11][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[11][6] ),
	.D(n280),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][5]  (
	.SI(\REG[11][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[11][5] ),
	.D(n279),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][4]  (
	.SI(\REG[11][3] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[11][4] ),
	.D(n278),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][3]  (
	.SI(\REG[11][2] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[11][3] ),
	.D(n277),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][2]  (
	.SI(\REG[11][1] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[11][2] ),
	.D(n276),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][1]  (
	.SI(\REG[11][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[11][1] ),
	.D(n275),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[11][0]  (
	.SI(\REG[10][7] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[11][0] ),
	.D(n274),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][7]  (
	.SI(\REG[7][6] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[7][7] ),
	.D(n249),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][6]  (
	.SI(\REG[7][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[7][6] ),
	.D(n248),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][5]  (
	.SI(\REG[7][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[7][5] ),
	.D(n247),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][4]  (
	.SI(\REG[7][3] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[7][4] ),
	.D(n246),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][3]  (
	.SI(\REG[7][2] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[7][3] ),
	.D(n245),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][2]  (
	.SI(\REG[7][1] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[7][2] ),
	.D(n244),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][1]  (
	.SI(\REG[7][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[7][1] ),
	.D(n243),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7][0]  (
	.SI(\REG[6][7] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[7][0] ),
	.D(n242),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][7]  (
	.SI(\REG[14][6] ),
	.SE(test_se),
	.RN(RST),
	.Q(\REG[14][7] ),
	.D(n305),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][6]  (
	.SI(\REG[14][5] ),
	.SE(test_se),
	.RN(RST),
	.Q(\REG[14][6] ),
	.D(n304),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][5]  (
	.SI(\REG[14][4] ),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(\REG[14][5] ),
	.D(n303),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][4]  (
	.SI(\REG[14][3] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[14][4] ),
	.D(n302),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][3]  (
	.SI(\REG[14][2] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[14][3] ),
	.D(n301),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][2]  (
	.SI(test_si3),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[14][2] ),
	.D(n300),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \REG_reg[14][1]  (
	.SI(\REG[14][0] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[14][1] ),
	.D(n299),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[14][0]  (
	.SI(\REG[13][7] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[14][0] ),
	.D(n298),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][7]  (
	.SI(\REG[10][6] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[10][7] ),
	.D(n273),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][6]  (
	.SI(\REG[10][5] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[10][6] ),
	.D(n272),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][5]  (
	.SI(\REG[10][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[10][5] ),
	.D(n271),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][4]  (
	.SI(\REG[10][3] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[10][4] ),
	.D(n270),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][3]  (
	.SI(\REG[10][2] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[10][3] ),
	.D(n269),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][2]  (
	.SI(\REG[10][1] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[10][2] ),
	.D(n268),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][1]  (
	.SI(\REG[10][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[10][1] ),
	.D(n267),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[10][0]  (
	.SI(\REG[9][7] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[10][0] ),
	.D(n266),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][7]  (
	.SI(\REG[6][6] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[6][7] ),
	.D(n241),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][6]  (
	.SI(\REG[6][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[6][6] ),
	.D(n240),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][5]  (
	.SI(\REG[6][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[6][5] ),
	.D(n239),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][4]  (
	.SI(\REG[6][3] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[6][4] ),
	.D(n238),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][3]  (
	.SI(\REG[6][2] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[6][3] ),
	.D(n237),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][2]  (
	.SI(\REG[6][1] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[6][2] ),
	.D(n236),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][1]  (
	.SI(\REG[6][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[6][1] ),
	.D(n235),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6][0]  (
	.SI(\REG[5][7] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[6][0] ),
	.D(n234),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][7]  (
	.SI(\REG[12][6] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][7] ),
	.D(n289),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][6]  (
	.SI(\REG[12][5] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][6] ),
	.D(n288),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][5]  (
	.SI(\REG[12][4] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][5] ),
	.D(n287),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][4]  (
	.SI(\REG[12][3] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][4] ),
	.D(n286),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][3]  (
	.SI(\REG[12][2] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][3] ),
	.D(n285),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][2]  (
	.SI(\REG[12][1] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][2] ),
	.D(n284),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][1]  (
	.SI(\REG[12][0] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][1] ),
	.D(n283),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[12][0]  (
	.SI(\REG[11][7] ),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[12][0] ),
	.D(n282),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][7]  (
	.SI(\REG[8][6] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[8][7] ),
	.D(n257),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][6]  (
	.SI(\REG[8][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][6] ),
	.D(n256),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][5]  (
	.SI(\REG[8][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][5] ),
	.D(n255),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][4]  (
	.SI(\REG[8][3] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][4] ),
	.D(n254),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][3]  (
	.SI(\REG[8][2] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][3] ),
	.D(n253),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][2]  (
	.SI(\REG[8][1] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][2] ),
	.D(n252),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][1]  (
	.SI(\REG[8][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][1] ),
	.D(n251),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[8][0]  (
	.SI(\REG[7][7] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[8][0] ),
	.D(n250),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][7]  (
	.SI(\REG[4][6] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[4][7] ),
	.D(n225),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][6]  (
	.SI(\REG[4][5] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[4][6] ),
	.D(n224),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][5]  (
	.SI(\REG[4][4] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(\REG[4][5] ),
	.D(n223),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][4]  (
	.SI(\REG[4][3] ),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[4][4] ),
	.D(n222),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][3]  (
	.SI(\REG[4][2] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[4][3] ),
	.D(n221),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][2]  (
	.SI(\REG[4][1] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[4][2] ),
	.D(n220),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][1]  (
	.SI(\REG[4][0] ),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[4][1] ),
	.D(n219),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4][0]  (
	.SI(REG_3[7]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(\REG[4][0] ),
	.D(n218),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][7]  (
	.SI(REG_0[6]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[7]),
	.D(n193),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][6]  (
	.SI(REG_0[5]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[6]),
	.D(n192),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][5]  (
	.SI(REG_0[4]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[5]),
	.D(n191),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][4]  (
	.SI(REG_0[3]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[4]),
	.D(n190),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][3]  (
	.SI(REG_0[2]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[3]),
	.D(n189),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][2]  (
	.SI(REG_0[1]),
	.SE(FE_OFN13_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[2]),
	.D(n188),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[7]  (
	.SI(RD_DATA[6]),
	.SE(test_se),
	.RN(RST),
	.Q(RD_DATA[7]),
	.D(n184),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[6]  (
	.SI(RD_DATA[5]),
	.SE(test_se),
	.RN(RST),
	.Q(RD_DATA[6]),
	.D(n183),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[5]  (
	.SI(RD_DATA[4]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA[5]),
	.D(n182),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[4]  (
	.SI(RD_DATA[3]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA[4]),
	.D(n181),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[3]  (
	.SI(RD_DATA[2]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA[3]),
	.D(n180),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[2]  (
	.SI(RD_DATA[1]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA[2]),
	.D(n179),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[1]  (
	.SI(RD_DATA[0]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA[1]),
	.D(n178),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_DATA_reg[0]  (
	.SI(RD_DATA_VALID),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA[0]),
	.D(n177),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][1]  (
	.SI(REG_2[0]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_2[1]),
	.D(n203),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][0]  (
	.SI(REG_2[7]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_3[0]),
	.D(n210),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][5]  (
	.SI(REG_1[4]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[5]),
	.D(n199),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][4]  (
	.SI(REG_1[3]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[4]),
	.D(n198),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][3]  (
	.SI(REG_1[2]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[3]),
	.D(n197),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][2]  (
	.SI(REG_1[1]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[2]),
	.D(n196),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][1]  (
	.SI(REG_1[0]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[1]),
	.D(n195),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][7]  (
	.SI(REG_1[6]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[7]),
	.D(n201),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][6]  (
	.SI(REG_1[5]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[6]),
	.D(n200),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1][0]  (
	.SI(REG_0[7]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_1[0]),
	.D(n194),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][1]  (
	.SI(REG_0[0]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN2_SYNC_REF_SCAN_RST),
	.Q(REG_0[1]),
	.D(n187),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \REG_reg[2][0]  (
	.SN(FE_OFN1_SYNC_REF_SCAN_RST),
	.SI(REG_1[7]),
	.SE(FE_OFN7_SE),
	.Q(REG_2[0]),
	.D(n202),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RD_DATA_VALID_reg (
	.SI(test_si1),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(RD_DATA_VALID),
	.D(n185),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][7]  (
	.SI(REG_3[6]),
	.SE(test_se),
	.RN(RST),
	.Q(REG_3[7]),
	.D(n217),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][6]  (
	.SI(REG_3[5]),
	.SE(test_se),
	.RN(RST),
	.Q(REG_3[6]),
	.D(n216),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][3]  (
	.SI(REG_3[2]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_3[3]),
	.D(n213),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][2]  (
	.SI(REG_3[1]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_3[2]),
	.D(n212),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \REG_reg[3][5]  (
	.SN(RST),
	.SI(REG_3[4]),
	.SE(test_se),
	.Q(REG_3[5]),
	.D(n215),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][4]  (
	.SI(REG_3[3]),
	.SE(test_se),
	.RN(RST),
	.Q(REG_3[4]),
	.D(n214),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3][1]  (
	.SI(REG_3[0]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(REG_3[1]),
	.D(n211),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][4]  (
	.SI(REG_2[3]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_2[4]),
	.D(n206),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \REG_reg[2][2]  (
	.SI(REG_2[1]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_2[2]),
	.D(n204),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \REG_reg[2][7]  (
	.SN(FE_OFN1_SYNC_REF_SCAN_RST),
	.SI(REG_2[6]),
	.SE(FE_OFN7_SE),
	.Q(REG_2[7]),
	.D(n209),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][5]  (
	.SI(REG_2[4]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_2[5]),
	.D(n207),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][6]  (
	.SI(REG_2[5]),
	.SE(FE_OFN7_SE),
	.RN(FE_OFN1_SYNC_REF_SCAN_RST),
	.Q(REG_2[6]),
	.D(n208),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2][3]  (
	.SI(test_si2),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_2[3]),
	.D(n205),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0][0]  (
	.SI(RD_DATA[7]),
	.SE(FE_OFN11_SE),
	.RN(FE_OFN0_SYNC_REF_SCAN_RST),
	.Q(REG_0[0]),
	.D(n186),
	.CK(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U140 (
	.Y(n169),
	.B(n340),
	.AN(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U141 (
	.Y(n155),
	.B(n340),
	.AN(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U142 (
	.Y(n160),
	.B(N12),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U143 (
	.Y(n163),
	.B(n341),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U144 (
	.Y(n157),
	.B(N13),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U145 (
	.Y(n152),
	.B(N13),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U146 (
	.Y(n338),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U147 (
	.Y(n336),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U148 (
	.Y(n339),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U150 (
	.Y(n361),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U152 (
	.Y(n153),
	.B(N11),
	.AN(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U153 (
	.Y(n167),
	.B(N11),
	.AN(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U154 (
	.Y(n166),
	.B(n152),
	.A(n167), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U155 (
	.Y(n168),
	.B(n152),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U156 (
	.Y(n170),
	.B(n157),
	.A(n167), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U157 (
	.Y(n171),
	.B(n157),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U158 (
	.Y(n156),
	.B(n153),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U159 (
	.Y(n158),
	.B(n155),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U160 (
	.Y(n172),
	.B(n160),
	.A(n167), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U161 (
	.Y(n173),
	.B(n160),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U162 (
	.Y(n174),
	.B(n163),
	.A(n167), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U163 (
	.Y(n176),
	.B(n163),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U164 (
	.Y(n150),
	.B(RD_EN),
	.AN(WR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U165 (
	.Y(n154),
	.B(n152),
	.A(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U166 (
	.Y(n159),
	.B(n153),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U167 (
	.Y(n161),
	.B(n155),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U168 (
	.Y(n162),
	.B(n153),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U169 (
	.Y(n165),
	.B(n155),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U170 (
	.Y(n151),
	.B(n153),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U171 (
	.Y(n149),
	.B(RD_EN),
	.AN(WR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U182 (
	.Y(n164),
	.B(N14),
	.AN(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U183 (
	.Y(n175),
	.B(n150),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U184 (
	.Y(n357),
	.A(WR_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U185 (
	.Y(n358),
	.A(WR_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U186 (
	.Y(n359),
	.A(WR_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U187 (
	.Y(n360),
	.A(WR_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U188 (
	.Y(n364),
	.A(WR_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U189 (
	.Y(n365),
	.A(WR_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U190 (
	.Y(n362),
	.A(WR_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U196 (
	.Y(n250),
	.B1(n166),
	.B0(n357),
	.A1N(n166),
	.A0N(\REG[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U197 (
	.Y(n251),
	.B1(n166),
	.B0(n358),
	.A1N(n166),
	.A0N(\REG[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U198 (
	.Y(n252),
	.B1(n166),
	.B0(n359),
	.A1N(n166),
	.A0N(\REG[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U199 (
	.Y(n253),
	.B1(n166),
	.B0(n360),
	.A1N(n166),
	.A0N(\REG[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U200 (
	.Y(n254),
	.B1(n166),
	.B0(n365),
	.A1N(n166),
	.A0N(\REG[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U201 (
	.Y(n255),
	.B1(n166),
	.B0(n364),
	.A1N(n166),
	.A0N(\REG[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U202 (
	.Y(n256),
	.B1(n166),
	.B0(n363),
	.A1N(n166),
	.A0N(\REG[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U203 (
	.Y(n257),
	.B1(n166),
	.B0(n362),
	.A1N(n166),
	.A0N(\REG[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U204 (
	.Y(n258),
	.B1(n168),
	.B0(n357),
	.A1N(n168),
	.A0N(\REG[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U205 (
	.Y(n259),
	.B1(n168),
	.B0(n358),
	.A1N(n168),
	.A0N(\REG[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U206 (
	.Y(n260),
	.B1(n168),
	.B0(n359),
	.A1N(n168),
	.A0N(\REG[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n261),
	.B1(n168),
	.B0(n360),
	.A1N(n168),
	.A0N(\REG[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n262),
	.B1(n168),
	.B0(n365),
	.A1N(n168),
	.A0N(\REG[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n263),
	.B1(n168),
	.B0(n364),
	.A1N(n168),
	.A0N(\REG[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n264),
	.B1(n168),
	.B0(n363),
	.A1N(n168),
	.A0N(\REG[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n265),
	.B1(n168),
	.B0(n362),
	.A1N(n168),
	.A0N(\REG[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n266),
	.B1(n170),
	.B0(n357),
	.A1N(n170),
	.A0N(\REG[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n267),
	.B1(n170),
	.B0(n358),
	.A1N(n170),
	.A0N(\REG[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n268),
	.B1(n170),
	.B0(n359),
	.A1N(n170),
	.A0N(\REG[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n269),
	.B1(n170),
	.B0(n360),
	.A1N(n170),
	.A0N(\REG[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n270),
	.B1(n170),
	.B0(n365),
	.A1N(n170),
	.A0N(\REG[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n271),
	.B1(n170),
	.B0(n364),
	.A1N(n170),
	.A0N(\REG[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n272),
	.B1(n170),
	.B0(n363),
	.A1N(n170),
	.A0N(\REG[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n273),
	.B1(n170),
	.B0(n362),
	.A1N(n170),
	.A0N(\REG[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n274),
	.B1(n171),
	.B0(n357),
	.A1N(n171),
	.A0N(\REG[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n275),
	.B1(n171),
	.B0(n358),
	.A1N(n171),
	.A0N(\REG[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n276),
	.B1(n171),
	.B0(n359),
	.A1N(n171),
	.A0N(\REG[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n277),
	.B1(n171),
	.B0(n360),
	.A1N(n171),
	.A0N(\REG[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n278),
	.B1(n171),
	.B0(n365),
	.A1N(n171),
	.A0N(\REG[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n279),
	.B1(n171),
	.B0(n364),
	.A1N(n171),
	.A0N(\REG[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n280),
	.B1(n171),
	.B0(n363),
	.A1N(n171),
	.A0N(\REG[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n281),
	.B1(n171),
	.B0(n362),
	.A1N(n171),
	.A0N(\REG[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n282),
	.B1(n172),
	.B0(n357),
	.A1N(n172),
	.A0N(\REG[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n283),
	.B1(n172),
	.B0(n358),
	.A1N(n172),
	.A0N(\REG[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n284),
	.B1(n172),
	.B0(n359),
	.A1N(n172),
	.A0N(\REG[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n285),
	.B1(n172),
	.B0(n360),
	.A1N(n172),
	.A0N(\REG[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n286),
	.B1(n172),
	.B0(n365),
	.A1N(n172),
	.A0N(\REG[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n287),
	.B1(n172),
	.B0(n364),
	.A1N(n172),
	.A0N(\REG[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n288),
	.B1(n172),
	.B0(n363),
	.A1N(n172),
	.A0N(\REG[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n289),
	.B1(n172),
	.B0(n362),
	.A1N(n172),
	.A0N(\REG[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n290),
	.B1(n173),
	.B0(n357),
	.A1N(n173),
	.A0N(\REG[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n291),
	.B1(n173),
	.B0(n358),
	.A1N(n173),
	.A0N(\REG[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U238 (
	.Y(n292),
	.B1(n173),
	.B0(n359),
	.A1N(n173),
	.A0N(\REG[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n293),
	.B1(n173),
	.B0(n360),
	.A1N(n173),
	.A0N(\REG[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U240 (
	.Y(n294),
	.B1(n173),
	.B0(n365),
	.A1N(n173),
	.A0N(\REG[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U241 (
	.Y(n295),
	.B1(n173),
	.B0(n364),
	.A1N(n173),
	.A0N(\REG[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U242 (
	.Y(n296),
	.B1(n173),
	.B0(n363),
	.A1N(n173),
	.A0N(\REG[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U243 (
	.Y(n297),
	.B1(n173),
	.B0(n362),
	.A1N(n173),
	.A0N(\REG[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U244 (
	.Y(n298),
	.B1(n174),
	.B0(n357),
	.A1N(n174),
	.A0N(\REG[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U245 (
	.Y(n299),
	.B1(n174),
	.B0(n358),
	.A1N(n174),
	.A0N(\REG[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U246 (
	.Y(n300),
	.B1(n174),
	.B0(n359),
	.A1N(n174),
	.A0N(\REG[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n301),
	.B1(n174),
	.B0(n360),
	.A1N(n174),
	.A0N(\REG[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U248 (
	.Y(n302),
	.B1(n174),
	.B0(n365),
	.A1N(n174),
	.A0N(\REG[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U249 (
	.Y(n303),
	.B1(n174),
	.B0(n364),
	.A1N(n174),
	.A0N(\REG[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U250 (
	.Y(n304),
	.B1(n174),
	.B0(n363),
	.A1N(n174),
	.A0N(\REG[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n305),
	.B1(n174),
	.B0(n362),
	.A1N(n174),
	.A0N(\REG[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U252 (
	.Y(n306),
	.B1(n176),
	.B0(n357),
	.A1N(n176),
	.A0N(\REG[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U253 (
	.Y(n307),
	.B1(n176),
	.B0(n358),
	.A1N(n176),
	.A0N(\REG[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U254 (
	.Y(n308),
	.B1(n176),
	.B0(n359),
	.A1N(n176),
	.A0N(\REG[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n309),
	.B1(n176),
	.B0(n360),
	.A1N(n176),
	.A0N(\REG[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U256 (
	.Y(n310),
	.B1(n176),
	.B0(n365),
	.A1N(n176),
	.A0N(\REG[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U257 (
	.Y(n311),
	.B1(n176),
	.B0(n364),
	.A1N(n176),
	.A0N(\REG[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U258 (
	.Y(n312),
	.B1(n176),
	.B0(n363),
	.A1N(n176),
	.A0N(\REG[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n313),
	.B1(n176),
	.B0(n362),
	.A1N(n176),
	.A0N(\REG[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U260 (
	.Y(n202),
	.B1(n156),
	.B0(n357),
	.A1N(n156),
	.A0N(REG_2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U261 (
	.Y(n209),
	.B1(n156),
	.B0(n362),
	.A1N(n156),
	.A0N(REG_2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U262 (
	.Y(n215),
	.B1(n158),
	.B0(n364),
	.A1N(n158),
	.A0N(REG_3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U263 (
	.Y(n177),
	.B1(n149),
	.B0(RD_DATA[0]),
	.A1(n361),
	.A0(N43), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U264 (
	.Y(N43),
	.S1(N13),
	.S0(N14),
	.D(n138),
	.C(n140),
	.B(n139),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U265 (
	.Y(n141),
	.S1(N12),
	.S0(N11),
	.D(REG_3[0]),
	.C(REG_2[0]),
	.B(REG_1[0]),
	.A(REG_0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U266 (
	.Y(n139),
	.S1(N12),
	.S0(N11),
	.D(\REG[11][0] ),
	.C(\REG[10][0] ),
	.B(\REG[9][0] ),
	.A(\REG[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U267 (
	.Y(n178),
	.B1(n149),
	.B0(RD_DATA[1]),
	.A1(n361),
	.A0(N42), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U268 (
	.Y(N42),
	.S1(N13),
	.S0(N14),
	.D(n142),
	.C(n144),
	.B(n143),
	.A(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U269 (
	.Y(n143),
	.S1(N12),
	.S0(N11),
	.D(\REG[11][1] ),
	.C(\REG[10][1] ),
	.B(\REG[9][1] ),
	.A(\REG[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U270 (
	.Y(n142),
	.S1(n336),
	.S0(n339),
	.D(\REG[15][1] ),
	.C(\REG[14][1] ),
	.B(\REG[13][1] ),
	.A(\REG[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U271 (
	.Y(n179),
	.B1(n149),
	.B0(RD_DATA[2]),
	.A1(n361),
	.A0(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U272 (
	.Y(N41),
	.S1(N13),
	.S0(N14),
	.D(n146),
	.C(n148),
	.B(n147),
	.A(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U273 (
	.Y(n314),
	.S1(n336),
	.S0(n338),
	.D(REG_3[2]),
	.C(REG_2[2]),
	.B(REG_1[2]),
	.A(REG_0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U274 (
	.Y(n147),
	.S1(n336),
	.S0(n338),
	.D(\REG[11][2] ),
	.C(\REG[10][2] ),
	.B(\REG[9][2] ),
	.A(\REG[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U275 (
	.Y(n180),
	.B1(n149),
	.B0(RD_DATA[3]),
	.A1(n361),
	.A0(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U276 (
	.Y(N40),
	.S1(N13),
	.S0(N14),
	.D(n315),
	.C(n317),
	.B(n316),
	.A(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U277 (
	.Y(n318),
	.S1(n336),
	.S0(n338),
	.D(REG_3[3]),
	.C(REG_2[3]),
	.B(REG_1[3]),
	.A(REG_0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U278 (
	.Y(n316),
	.S1(n336),
	.S0(n338),
	.D(\REG[11][3] ),
	.C(\REG[10][3] ),
	.B(\REG[9][3] ),
	.A(\REG[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U279 (
	.Y(n181),
	.B1(n149),
	.B0(RD_DATA[4]),
	.A1(n361),
	.A0(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U280 (
	.Y(N39),
	.S1(N13),
	.S0(N14),
	.D(n319),
	.C(n321),
	.B(n320),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U281 (
	.Y(n322),
	.S1(n336),
	.S0(n339),
	.D(REG_3[4]),
	.C(REG_2[4]),
	.B(REG_1[4]),
	.A(REG_0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U282 (
	.Y(n320),
	.S1(n336),
	.S0(n338),
	.D(\REG[11][4] ),
	.C(\REG[10][4] ),
	.B(\REG[9][4] ),
	.A(\REG[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U283 (
	.Y(n182),
	.B1(n149),
	.B0(RD_DATA[5]),
	.A1(n361),
	.A0(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U284 (
	.Y(N38),
	.S1(N13),
	.S0(N14),
	.D(n323),
	.C(n325),
	.B(n324),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U285 (
	.Y(n326),
	.S1(N12),
	.S0(n339),
	.D(REG_3[5]),
	.C(REG_2[5]),
	.B(REG_1[5]),
	.A(REG_0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U286 (
	.Y(n324),
	.S1(N12),
	.S0(n339),
	.D(\REG[11][5] ),
	.C(\REG[10][5] ),
	.B(\REG[9][5] ),
	.A(\REG[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U287 (
	.Y(n183),
	.B1(n149),
	.B0(RD_DATA[6]),
	.A1(n361),
	.A0(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U288 (
	.Y(N37),
	.S1(N13),
	.S0(N14),
	.D(n327),
	.C(n329),
	.B(n328),
	.A(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U289 (
	.Y(n330),
	.S1(N12),
	.S0(n339),
	.D(REG_3[6]),
	.C(REG_2[6]),
	.B(REG_1[6]),
	.A(REG_0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U290 (
	.Y(n328),
	.S1(N12),
	.S0(n339),
	.D(\REG[11][6] ),
	.C(\REG[10][6] ),
	.B(\REG[9][6] ),
	.A(\REG[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U291 (
	.Y(n184),
	.B1(n149),
	.B0(RD_DATA[7]),
	.A1(n361),
	.A0(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U292 (
	.Y(N36),
	.S1(N13),
	.S0(N14),
	.D(n331),
	.C(n333),
	.B(n332),
	.A(n334), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U293 (
	.Y(n334),
	.S1(N12),
	.S0(n339),
	.D(REG_3[7]),
	.C(REG_2[7]),
	.B(REG_1[7]),
	.A(REG_0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U294 (
	.Y(n332),
	.S1(N12),
	.S0(n339),
	.D(\REG[11][7] ),
	.C(\REG[10][7] ),
	.B(\REG[9][7] ),
	.A(\REG[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U295 (
	.Y(n145),
	.S1(N12),
	.S0(n338),
	.D(REG_3[1]),
	.C(REG_2[1]),
	.B(REG_1[1]),
	.A(REG_0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U296 (
	.Y(n140),
	.S1(N12),
	.S0(N11),
	.D(\REG[7][0] ),
	.C(\REG[6][0] ),
	.B(\REG[5][0] ),
	.A(\REG[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U297 (
	.Y(n144),
	.S1(N12),
	.S0(n338),
	.D(\REG[7][1] ),
	.C(\REG[6][1] ),
	.B(\REG[5][1] ),
	.A(\REG[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U298 (
	.Y(n148),
	.S1(n336),
	.S0(n338),
	.D(\REG[7][2] ),
	.C(\REG[6][2] ),
	.B(\REG[5][2] ),
	.A(\REG[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U299 (
	.Y(n317),
	.S1(n336),
	.S0(n338),
	.D(\REG[7][3] ),
	.C(\REG[6][3] ),
	.B(\REG[5][3] ),
	.A(\REG[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U300 (
	.Y(n321),
	.S1(n336),
	.S0(n338),
	.D(\REG[7][4] ),
	.C(\REG[6][4] ),
	.B(\REG[5][4] ),
	.A(\REG[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U301 (
	.Y(n325),
	.S1(N12),
	.S0(n339),
	.D(\REG[7][5] ),
	.C(\REG[6][5] ),
	.B(\REG[5][5] ),
	.A(\REG[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U302 (
	.Y(n329),
	.S1(N12),
	.S0(n339),
	.D(\REG[7][6] ),
	.C(\REG[6][6] ),
	.B(\REG[5][6] ),
	.A(\REG[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U303 (
	.Y(n333),
	.S1(N12),
	.S0(n339),
	.D(\REG[7][7] ),
	.C(\REG[6][7] ),
	.B(\REG[5][7] ),
	.A(\REG[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U304 (
	.Y(n138),
	.S1(n336),
	.S0(n338),
	.D(\REG[15][0] ),
	.C(\REG[14][0] ),
	.B(\REG[13][0] ),
	.A(\REG[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U305 (
	.Y(n146),
	.S1(n336),
	.S0(n338),
	.D(\REG[15][2] ),
	.C(\REG[14][2] ),
	.B(\REG[13][2] ),
	.A(\REG[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U306 (
	.Y(n315),
	.S1(n336),
	.S0(n338),
	.D(\REG[15][3] ),
	.C(\REG[14][3] ),
	.B(\REG[13][3] ),
	.A(\REG[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U307 (
	.Y(n319),
	.S1(n336),
	.S0(n338),
	.D(\REG[15][4] ),
	.C(\REG[14][4] ),
	.B(\REG[13][4] ),
	.A(\REG[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U308 (
	.Y(n323),
	.S1(N12),
	.S0(n339),
	.D(\REG[15][5] ),
	.C(\REG[14][5] ),
	.B(\REG[13][5] ),
	.A(\REG[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U309 (
	.Y(n327),
	.S1(N12),
	.S0(n339),
	.D(\REG[15][6] ),
	.C(\REG[14][6] ),
	.B(\REG[13][6] ),
	.A(\REG[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U310 (
	.Y(n331),
	.S1(N12),
	.S0(n339),
	.D(\REG[15][7] ),
	.C(\REG[14][7] ),
	.B(\REG[13][7] ),
	.A(\REG[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U311 (
	.Y(n340),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U312 (
	.Y(n363),
	.A(WR_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U313 (
	.Y(n186),
	.B1(n357),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U314 (
	.Y(n187),
	.B1(n358),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U315 (
	.Y(n188),
	.B1(n359),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U316 (
	.Y(n189),
	.B1(n360),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U317 (
	.Y(n190),
	.B1(n365),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U318 (
	.Y(n191),
	.B1(n364),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U319 (
	.Y(n192),
	.B1(n363),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U320 (
	.Y(n193),
	.B1(n362),
	.B0(n151),
	.A1N(n151),
	.A0N(REG_0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U321 (
	.Y(n194),
	.B1(n154),
	.B0(n357),
	.A1N(n154),
	.A0N(REG_1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U322 (
	.Y(n195),
	.B1(n154),
	.B0(n358),
	.A1N(n154),
	.A0N(REG_1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U323 (
	.Y(n196),
	.B1(n154),
	.B0(n359),
	.A1N(n154),
	.A0N(REG_1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U324 (
	.Y(n197),
	.B1(n154),
	.B0(n360),
	.A1N(n154),
	.A0N(REG_1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U325 (
	.Y(n198),
	.B1(n154),
	.B0(n365),
	.A1N(n154),
	.A0N(REG_1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U326 (
	.Y(n199),
	.B1(n154),
	.B0(n364),
	.A1N(n154),
	.A0N(REG_1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U327 (
	.Y(n200),
	.B1(n154),
	.B0(n363),
	.A1N(n154),
	.A0N(REG_1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U328 (
	.Y(n201),
	.B1(n154),
	.B0(n362),
	.A1N(n154),
	.A0N(REG_1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U329 (
	.Y(n218),
	.B1(n159),
	.B0(n357),
	.A1N(n159),
	.A0N(\REG[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U330 (
	.Y(n219),
	.B1(n159),
	.B0(n358),
	.A1N(n159),
	.A0N(\REG[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U331 (
	.Y(n220),
	.B1(n159),
	.B0(n359),
	.A1N(n159),
	.A0N(\REG[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U332 (
	.Y(n221),
	.B1(n159),
	.B0(n360),
	.A1N(n159),
	.A0N(\REG[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U333 (
	.Y(n222),
	.B1(n159),
	.B0(n365),
	.A1N(n159),
	.A0N(\REG[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U334 (
	.Y(n223),
	.B1(n159),
	.B0(n364),
	.A1N(n159),
	.A0N(\REG[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U335 (
	.Y(n224),
	.B1(n159),
	.B0(n363),
	.A1N(n159),
	.A0N(\REG[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U336 (
	.Y(n225),
	.B1(n159),
	.B0(n362),
	.A1N(n159),
	.A0N(\REG[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U337 (
	.Y(n226),
	.B1(n161),
	.B0(n357),
	.A1N(n161),
	.A0N(\REG[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U338 (
	.Y(n227),
	.B1(n161),
	.B0(n358),
	.A1N(n161),
	.A0N(\REG[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U339 (
	.Y(n228),
	.B1(n161),
	.B0(n359),
	.A1N(n161),
	.A0N(\REG[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U340 (
	.Y(n229),
	.B1(n161),
	.B0(n360),
	.A1N(n161),
	.A0N(\REG[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U341 (
	.Y(n230),
	.B1(n161),
	.B0(n365),
	.A1N(n161),
	.A0N(\REG[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U342 (
	.Y(n231),
	.B1(n161),
	.B0(n364),
	.A1N(n161),
	.A0N(\REG[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U343 (
	.Y(n232),
	.B1(n161),
	.B0(n363),
	.A1N(n161),
	.A0N(\REG[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U344 (
	.Y(n233),
	.B1(n161),
	.B0(n362),
	.A1N(n161),
	.A0N(\REG[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U345 (
	.Y(n234),
	.B1(n162),
	.B0(n357),
	.A1N(n162),
	.A0N(\REG[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U346 (
	.Y(n235),
	.B1(n162),
	.B0(n358),
	.A1N(n162),
	.A0N(\REG[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U347 (
	.Y(n236),
	.B1(n162),
	.B0(n359),
	.A1N(n162),
	.A0N(\REG[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U348 (
	.Y(n237),
	.B1(n162),
	.B0(n360),
	.A1N(n162),
	.A0N(\REG[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U349 (
	.Y(n238),
	.B1(n162),
	.B0(n365),
	.A1N(n162),
	.A0N(\REG[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U350 (
	.Y(n239),
	.B1(n162),
	.B0(n364),
	.A1N(n162),
	.A0N(\REG[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U351 (
	.Y(n240),
	.B1(n162),
	.B0(n363),
	.A1N(n162),
	.A0N(\REG[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U352 (
	.Y(n241),
	.B1(n162),
	.B0(n362),
	.A1N(n162),
	.A0N(\REG[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U353 (
	.Y(n242),
	.B1(n165),
	.B0(n357),
	.A1N(n165),
	.A0N(\REG[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U354 (
	.Y(n243),
	.B1(n165),
	.B0(n358),
	.A1N(n165),
	.A0N(\REG[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U355 (
	.Y(n244),
	.B1(n165),
	.B0(n359),
	.A1N(n165),
	.A0N(\REG[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U356 (
	.Y(n245),
	.B1(n165),
	.B0(n360),
	.A1N(n165),
	.A0N(\REG[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U357 (
	.Y(n246),
	.B1(n165),
	.B0(n365),
	.A1N(n165),
	.A0N(\REG[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U358 (
	.Y(n247),
	.B1(n165),
	.B0(n364),
	.A1N(n165),
	.A0N(\REG[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U359 (
	.Y(n248),
	.B1(n165),
	.B0(n363),
	.A1N(n165),
	.A0N(\REG[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U360 (
	.Y(n249),
	.B1(n165),
	.B0(n362),
	.A1N(n165),
	.A0N(\REG[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U361 (
	.Y(n203),
	.B1(n156),
	.B0(n358),
	.A1N(n156),
	.A0N(REG_2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U362 (
	.Y(n204),
	.B1(n156),
	.B0(n359),
	.A1N(n156),
	.A0N(REG_2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U363 (
	.Y(n205),
	.B1(n156),
	.B0(n360),
	.A1N(n156),
	.A0N(REG_2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U364 (
	.Y(n206),
	.B1(n156),
	.B0(n365),
	.A1N(n156),
	.A0N(REG_2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U365 (
	.Y(n207),
	.B1(n156),
	.B0(n364),
	.A1N(n156),
	.A0N(REG_2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U366 (
	.Y(n208),
	.B1(n156),
	.B0(n363),
	.A1N(n156),
	.A0N(REG_2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U367 (
	.Y(n210),
	.B1(n158),
	.B0(n357),
	.A1N(n158),
	.A0N(REG_3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U368 (
	.Y(n211),
	.B1(n158),
	.B0(n358),
	.A1N(n158),
	.A0N(REG_3[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U369 (
	.Y(n212),
	.B1(n158),
	.B0(n359),
	.A1N(n158),
	.A0N(REG_3[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U370 (
	.Y(n213),
	.B1(n158),
	.B0(n360),
	.A1N(n158),
	.A0N(REG_3[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U371 (
	.Y(n214),
	.B1(n158),
	.B0(n365),
	.A1N(n158),
	.A0N(REG_3[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U372 (
	.Y(n216),
	.B1(n158),
	.B0(n363),
	.A1N(n158),
	.A0N(REG_3[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U373 (
	.Y(n217),
	.B1(n158),
	.B0(n362),
	.A1N(n158),
	.A0N(REG_3[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U374 (
	.Y(n185),
	.B0(n149),
	.A1N(n150),
	.A0N(RD_DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U375 (
	.Y(n341),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_GATE (
	CLK, 
	CLK_EN, 
	GATED_CLK, 
	VDD, 
	VSS);
   input CLK;
   input CLK_EN;
   output GATED_CLK;
   inout VDD;
   inout VSS;

   // Module instantiations
   TLATNCAX12M U0_TLATNCAX12M (
	.ECK(GATED_CLK),
	.E(CLK_EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPERAND_WIDTH8_FUN_WIDTH4_test_1 (
	CLK, 
	RST, 
	A, 
	B, 
	ALU_FUN, 
	ALU_EN, 
	ALU_OUT, 
	OUT_VALID, 
	test_si, 
	test_se, 
	FE_OFN7_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input ALU_EN;
   output [15:0] ALU_OUT;
   output OUT_VALID;
   input test_si;
   input test_se;
   input FE_OFN7_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N88;
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N154;
   wire N155;
   wire N157;
   wire N158;
   wire N159;
   wire N160;
   wire N161;
   wire N162;
   wire N163;
   wire N164;
   wire N165;
   wire N166;
   wire N167;
   wire N168;
   wire N169;
   wire N170;
   wire N171;
   wire N172;
   wire N173;
   wire \U3/U1/Z_0 ;
   wire \U3/U1/Z_1 ;
   wire \U3/U1/Z_4 ;
   wire \U3/U1/Z_6 ;
   wire \U3/U1/Z_7 ;
   wire \U3/U2/Z_0 ;
   wire \U3/U2/Z_1 ;
   wire \U3/U2/Z_2 ;
   wire \U3/U2/Z_3 ;
   wire \U3/U2/Z_4 ;
   wire \U3/U2/Z_5 ;
   wire \U3/U2/Z_6 ;
   wire \U3/U2/Z_7 ;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n3;
   wire n4;
   wire n5;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;

   // Module instantiations
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[15]),
	.D(N172),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[14]),
	.D(N171),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[13]),
	.D(N170),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[12]),
	.D(N169),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[11]),
	.D(N168),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[10]),
	.D(N167),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[9]),
	.D(N166),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[8]),
	.D(N165),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[7]),
	.D(N164),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[6]),
	.D(N163),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[5]),
	.D(N162),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[4]),
	.D(N161),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[3]),
	.D(N160),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[2]),
	.D(N159),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[1]),
	.D(N158),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN7_SE),
	.RN(RST),
	.Q(ALU_OUT[0]),
	.D(N157),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M OUT_VALID_reg (
	.SI(ALU_OUT[15]),
	.SE(test_se),
	.RN(RST),
	.Q(OUT_VALID),
	.D(N173),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U23 (
	.Y(n68),
	.B(n70),
	.AN(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U24 (
	.Y(n93),
	.B(n142),
	.A(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n150),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n151),
	.A(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n147),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n148),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U31 (
	.Y(n72),
	.B0(n142),
	.A1N(n130),
	.A0N(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U32 (
	.Y(n140),
	.B(n149),
	.A(n154), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U33 (
	.Y(n82),
	.B(n144),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U34 (
	.Y(n83),
	.B(n131),
	.A(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U35 (
	.Y(n130),
	.B(n152),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U36 (
	.Y(n77),
	.B(n139),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U37 (
	.Y(n81),
	.B(n145),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U38 (
	.Y(n80),
	.B(n143),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U39 (
	.Y(n86),
	.B(n131),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U40 (
	.Y(n79),
	.B(n143),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U41 (
	.Y(n142),
	.B(n140),
	.A(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U42 (
	.Y(n75),
	.B(n139),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U43 (
	.Y(n132),
	.B(n140),
	.A(n139), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BBX1M U44 (
	.Y(N173),
	.D(n74),
	.C(n73),
	.BN(n72),
	.AN(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U45 (
	.Y(n73),
	.C(n83),
	.B(n82),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U46 (
	.Y(n74),
	.D(n78),
	.C(n77),
	.B(n76),
	.AN(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U47 (
	.Y(n76),
	.C(n81),
	.B(n80),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U48 (
	.Y(n78),
	.B(n145),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U49 (
	.Y(n67),
	.B(n131),
	.A(n139), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U50 (
	.Y(n69),
	.B(n140),
	.A(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U51 (
	.Y(n70),
	.B(n145),
	.A(n131), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U52 (
	.Y(n143),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U53 (
	.Y(n144),
	.B(ALU_FUN[0]),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U54 (
	.Y(n139),
	.B(ALU_FUN[1]),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U55 (
	.Y(n145),
	.B(ALU_FUN[2]),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U56 (
	.Y(n131),
	.B(ALU_FUN[0]),
	.A(n154), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U57 (
	.Y(n50),
	.A(\U3/U2/Z_6 ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U58 (
	.Y(n141),
	.B(ALU_FUN[3]),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U59 (
	.Y(N166),
	.B0(n84),
	.A1N(n151),
	.A0N(N115), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U60 (
	.Y(N167),
	.B0(n84),
	.A1N(n151),
	.A0N(N116), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U61 (
	.Y(N168),
	.B0(n84),
	.A1N(n151),
	.A0N(N117), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U62 (
	.Y(N169),
	.B0(n84),
	.A1N(n151),
	.A0N(N118), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U63 (
	.Y(N170),
	.B0(n84),
	.A1N(n151),
	.A0N(N119), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U64 (
	.Y(N171),
	.B0(n84),
	.A1N(n151),
	.A0N(N120), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U65 (
	.Y(N172),
	.B0(n84),
	.A1N(n151),
	.A0N(N121), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U66 (
	.Y(n71),
	.B0(n146),
	.A1N(n70),
	.A0N(N154), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U67 (
	.Y(n146),
	.B0(N155),
	.A1N(n69),
	.A0N(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U68 (
	.Y(n153),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U69 (
	.Y(n154),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U70 (
	.Y(n149),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U71 (
	.Y(n152),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U72 (
	.Y(n49),
	.A(\U3/U2/Z_4 ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U73 (
	.Y(n84),
	.C0(n72),
	.B0(n82),
	.A1(n147),
	.A0(N105), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U74 (
	.Y(\U3/U2/Z_4 ),
	.B1(n54),
	.B0(n68),
	.A1(n62),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U75 (
	.Y(\U3/U2/Z_6 ),
	.B1(n52),
	.B0(n68),
	.A1(n60),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U76 (
	.Y(\U3/U2/Z_5 ),
	.B1(n53),
	.B0(n68),
	.A1(n61),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U77 (
	.Y(\U3/U2/Z_2 ),
	.B1(n56),
	.B0(n68),
	.A1(n64),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U78 (
	.Y(\U3/U2/Z_3 ),
	.B1(n55),
	.B0(n68),
	.A1(n63),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U79 (
	.Y(\U3/U1/Z_1 ),
	.B1(n65),
	.B0(n68),
	.A1(n57),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U80 (
	.Y(\U3/U2/Z_1 ),
	.B1(n57),
	.B0(n68),
	.A1(n65),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U81 (
	.Y(\U3/U1/Z_4 ),
	.B1(n62),
	.B0(n68),
	.A1(n54),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U82 (
	.Y(\U3/U1/Z_6 ),
	.B1(n60),
	.B0(n68),
	.A1(n52),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U83 (
	.Y(\U3/U2/Z_7 ),
	.B1(n51),
	.B0(n68),
	.A1(n59),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U84 (
	.Y(\U3/U1/Z_7 ),
	.B1(n59),
	.B0(n68),
	.A1(n67),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U85 (
	.Y(\U3/U2/Z_0 ),
	.B1(n58),
	.B0(n68),
	.A1(n66),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U86 (
	.Y(\U3/U1/Z_0 ),
	.B1(n66),
	.B0(n68),
	.A1(n58),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U87 (
	.Y(N165),
	.C0(n85),
	.B0(n84),
	.A1N(N96),
	.A0(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U88 (
	.Y(n85),
	.B1(n151),
	.B0(N114),
	.A1N(n59),
	.A0N(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U89 (
	.Y(N159),
	.C(n120),
	.B(n119),
	.A(n118), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U90 (
	.Y(n118),
	.B1(n150),
	.B0(N90),
	.A1(n147),
	.A0(N99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U91 (
	.Y(n120),
	.C0(n121),
	.B1(n64),
	.B0(n82),
	.A1(A[3]),
	.A0(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U92 (
	.Y(n119),
	.C1(n78),
	.C0(N124),
	.B1(A[2]),
	.B0(n77),
	.A1(n151),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U93 (
	.Y(N160),
	.C(n114),
	.B(n113),
	.A(n112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U94 (
	.Y(n112),
	.B1(n150),
	.B0(N91),
	.A1(n147),
	.A0(N100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U95 (
	.Y(n114),
	.C0(n115),
	.B1(n63),
	.B0(n82),
	.A1(A[4]),
	.A0(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U96 (
	.Y(n113),
	.C1(n78),
	.C0(N125),
	.B1(A[3]),
	.B0(n77),
	.A1(n151),
	.A0(N109), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U97 (
	.Y(N161),
	.C(n108),
	.B(n107),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U98 (
	.Y(n106),
	.B1(n150),
	.B0(N92),
	.A1(n147),
	.A0(N101), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U99 (
	.Y(n108),
	.C0(n109),
	.B1(n62),
	.B0(n82),
	.A1(A[5]),
	.A0(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U100 (
	.Y(n107),
	.C1(n78),
	.C0(N126),
	.B1(A[4]),
	.B0(n77),
	.A1(n151),
	.A0(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U101 (
	.Y(N162),
	.C(n102),
	.B(n101),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U102 (
	.Y(n100),
	.B1(n150),
	.B0(N93),
	.A1(n147),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U103 (
	.Y(n102),
	.C0(n103),
	.B1(n61),
	.B0(n82),
	.A1(A[6]),
	.A0(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U104 (
	.Y(n101),
	.C1(n78),
	.C0(N127),
	.B1(A[5]),
	.B0(n77),
	.A1(n151),
	.A0(N111), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U105 (
	.Y(N163),
	.C(n96),
	.B(n95),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U106 (
	.Y(n94),
	.B1(n150),
	.B0(N94),
	.A1(n147),
	.A0(N103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U107 (
	.Y(n96),
	.C0(n97),
	.B1(n60),
	.B0(n82),
	.A1(A[7]),
	.A0(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U108 (
	.Y(n95),
	.C1(n78),
	.C0(N128),
	.B1(A[6]),
	.B0(n77),
	.A1(n151),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U109 (
	.Y(N164),
	.C(n89),
	.B(n88),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U110 (
	.Y(n88),
	.B1(n151),
	.B0(N113),
	.A1(n78),
	.A0(N129), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U111 (
	.Y(n87),
	.B1(n150),
	.B0(N95),
	.A1(n147),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U112 (
	.Y(n89),
	.C0(n90),
	.B1(A[7]),
	.B0(n77),
	.A1(n59),
	.A0(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U113 (
	.Y(n64),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U114 (
	.Y(n63),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U115 (
	.Y(n62),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U116 (
	.Y(n61),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U117 (
	.Y(n60),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U118 (
	.Y(n59),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA22X2M U119 (
	.Y(n3),
	.B1(n64),
	.B0(n68),
	.A1(n56),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OA22X2M U120 (
	.Y(n4),
	.B1(n63),
	.B0(n68),
	.A1(n55),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OA22X2M U121 (
	.Y(n5),
	.B1(n61),
	.B0(n68),
	.A1(n53),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U122 (
	.Y(n136),
	.C1(n132),
	.C0(n65),
	.B1(n138),
	.B0(B[0]),
	.A1(n58),
	.A0(n137), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U123 (
	.Y(n138),
	.C0(n82),
	.B1(n66),
	.B0(n72),
	.A1(A[0]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U124 (
	.Y(n137),
	.C0(n77),
	.B1(n93),
	.B0(A[0]),
	.A1(n66),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U125 (
	.Y(n127),
	.C1(n86),
	.C0(n66),
	.B1(n129),
	.B0(B[1]),
	.A1(n57),
	.A0(n128), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U126 (
	.Y(n129),
	.C0(n82),
	.B1(n65),
	.B0(n72),
	.A1(A[1]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U127 (
	.Y(n128),
	.C0(n77),
	.B1(n93),
	.B0(A[1]),
	.A1(n65),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U128 (
	.Y(n121),
	.C1(n86),
	.C0(n65),
	.B1(n123),
	.B0(B[2]),
	.A1(n56),
	.A0(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U129 (
	.Y(n123),
	.C0(n82),
	.B1(n64),
	.B0(n72),
	.A1(A[2]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U130 (
	.Y(n122),
	.C0(n77),
	.B1(n93),
	.B0(A[2]),
	.A1(n64),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U131 (
	.Y(n115),
	.C1(n86),
	.C0(n64),
	.B1(n117),
	.B0(B[3]),
	.A1(n55),
	.A0(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U132 (
	.Y(n117),
	.C0(n82),
	.B1(n63),
	.B0(n72),
	.A1(A[3]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U133 (
	.Y(n116),
	.C0(n77),
	.B1(n93),
	.B0(A[3]),
	.A1(n63),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U134 (
	.Y(n109),
	.C1(n86),
	.C0(n63),
	.B1(n111),
	.B0(B[4]),
	.A1(n54),
	.A0(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U135 (
	.Y(n111),
	.C0(n82),
	.B1(n62),
	.B0(n72),
	.A1(A[4]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U136 (
	.Y(n110),
	.C0(n77),
	.B1(n93),
	.B0(A[4]),
	.A1(n62),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U137 (
	.Y(n103),
	.C1(n86),
	.C0(n62),
	.B1(n105),
	.B0(B[5]),
	.A1(n53),
	.A0(n104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U138 (
	.Y(n105),
	.C0(n82),
	.B1(n61),
	.B0(n72),
	.A1(A[5]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U139 (
	.Y(n104),
	.C0(n77),
	.B1(n93),
	.B0(A[5]),
	.A1(n61),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U140 (
	.Y(n97),
	.C1(n86),
	.C0(n61),
	.B1(n99),
	.B0(B[6]),
	.A1(n52),
	.A0(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U141 (
	.Y(n99),
	.C0(n82),
	.B1(n60),
	.B0(n72),
	.A1(A[6]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U142 (
	.Y(n98),
	.C0(n77),
	.B1(n93),
	.B0(A[6]),
	.A1(n60),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U143 (
	.Y(n90),
	.C1(n86),
	.C0(n60),
	.B1(n92),
	.B0(B[7]),
	.A1(n51),
	.A0(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U144 (
	.Y(n92),
	.C0(n82),
	.B1(n59),
	.B0(n72),
	.A1(A[7]),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U145 (
	.Y(n91),
	.C0(n77),
	.B1(n93),
	.B0(A[7]),
	.A1(n59),
	.A0(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U146 (
	.Y(n65),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U147 (
	.Y(n66),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U148 (
	.Y(N158),
	.C(n126),
	.B(n125),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U149 (
	.Y(n124),
	.B1(n150),
	.B0(N89),
	.A1(n147),
	.A0(N98), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U150 (
	.Y(n126),
	.C0(n127),
	.B1(n65),
	.B0(n82),
	.A1(A[2]),
	.A0(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U151 (
	.Y(n125),
	.C1(n78),
	.C0(N123),
	.B1(A[1]),
	.B0(n77),
	.A1(n151),
	.A0(N107), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U152 (
	.Y(N157),
	.C(n135),
	.B(n134),
	.A(n133), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U153 (
	.Y(n133),
	.B0(n71),
	.A1(n150),
	.A0(N88), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U154 (
	.Y(n135),
	.C0(n136),
	.B1(A[0]),
	.B0(n77),
	.A1(n66),
	.A0(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U155 (
	.Y(n134),
	.C1(n151),
	.C0(N106),
	.B1(n78),
	.B0(N122),
	.A1(n147),
	.A0(N97), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U162 (
	.Y(n58),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U163 (
	.Y(n51),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U164 (
	.Y(n52),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U165 (
	.Y(n56),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U166 (
	.Y(n57),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U167 (
	.Y(n55),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U168 (
	.Y(n54),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U169 (
	.Y(n53),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U170 (
	.Y(n15),
	.B(\U3/U1/Z_0 ),
	.AN(\U3/U2/Z_0 ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U171 (
	.Y(n16),
	.B1(n15),
	.B0(\U3/U2/Z_1 ),
	.A1N(\U3/U1/Z_1 ),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U172 (
	.Y(n44),
	.B(\U3/U2/Z_6 ),
	.AN(\U3/U1/Z_6 ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U173 (
	.Y(n43),
	.B(n5),
	.A(\U3/U2/Z_5 ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U174 (
	.Y(n23),
	.B(\U3/U2/Z_4 ),
	.AN(\U3/U1/Z_4 ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U175 (
	.Y(n48),
	.D(n23),
	.C(n43),
	.B(n44),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U176 (
	.Y(n22),
	.B(n4),
	.A(\U3/U2/Z_3 ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U177 (
	.Y(n17),
	.B(n3),
	.A(\U3/U2/Z_2 ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U178 (
	.Y(n47),
	.B(n17),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U179 (
	.Y(n46),
	.B(\U3/U1/Z_7 ),
	.AN(\U3/U2/Z_7 ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U180 (
	.Y(n19),
	.B(\U3/U2/Z_0 ),
	.AN(\U3/U1/Z_0 ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U181 (
	.Y(n18),
	.B0(\U3/U2/Z_1 ),
	.A1N(\U3/U1/Z_1 ),
	.A0N(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U182 (
	.Y(n20),
	.C0(n17),
	.B0(n18),
	.A1(n19),
	.A0(\U3/U1/Z_1 ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U183 (
	.Y(n21),
	.C0(n20),
	.B1(n4),
	.B0(\U3/U2/Z_3 ),
	.A1(n3),
	.A0(\U3/U2/Z_2 ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U184 (
	.Y(n24),
	.B1(n49),
	.B0(\U3/U1/Z_4 ),
	.A2(n21),
	.A1(n22),
	.A0(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U185 (
	.Y(n25),
	.B0(n24),
	.A1(n5),
	.A0(\U3/U2/Z_5 ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U186 (
	.Y(n45),
	.B1(n50),
	.B0(\U3/U1/Z_6 ),
	.A2(n25),
	.A1(n43),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U187 (
	.Y(N155),
	.B1(n45),
	.B0(n46),
	.A1N(\U3/U1/Z_7 ),
	.A0(\U3/U2/Z_7 ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U188 (
	.Y(N154),
	.D(n46),
	.C(N155),
	.B(n47),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW_div_uns_0 div_48 (
	.a({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.b({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.quotient({ N129,
		N128,
		N127,
		N126,
		N125,
		N124,
		N123,
		N122 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW01_sub_0 sub_36 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.DIFF({ N105,
		N104,
		N103,
		N102,
		N101,
		N100,
		N99,
		N98,
		N97 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW01_add_0 add_30 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.SUM({ N96,
		N95,
		N94,
		N93,
		N92,
		N91,
		N90,
		N89,
		N88 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW02_mult_0 mult_42 (
	.A({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.TC(1'b0),
	.PRODUCT({ N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109,
		N108,
		N107,
		N106 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[1][4] ;
   wire \u_div/CryTmp[1][5] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][4] ;
   wire \u_div/CryTmp[2][5] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[3][4] ;
   wire \u_div/CryTmp[3][5] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[4][4] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[6][2] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;

   // Module instantiations
   ADDFX2M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/CryTmp[0][1] ),
	.B(n17),
	.A(\u_div/PartRem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_1  (
	.S(\u_div/SumTmp[1][1] ),
	.CO(\u_div/CryTmp[1][2] ),
	.CI(\u_div/CryTmp[1][1] ),
	.B(n17),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_6  (
	.S(\u_div/SumTmp[1][6] ),
	.CO(\u_div/CryTmp[1][7] ),
	.CI(\u_div/CryTmp[1][6] ),
	.B(n12),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_5  (
	.S(\u_div/SumTmp[2][5] ),
	.CO(\u_div/CryTmp[2][6] ),
	.CI(\u_div/CryTmp[2][5] ),
	.B(n13),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_3  (
	.S(\u_div/SumTmp[4][3] ),
	.CO(\u_div/CryTmp[4][4] ),
	.CI(\u_div/CryTmp[4][3] ),
	.B(n15),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_2  (
	.S(\u_div/SumTmp[5][2] ),
	.CO(\u_div/CryTmp[5][3] ),
	.CI(\u_div/CryTmp[5][2] ),
	.B(n16),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_6_1  (
	.S(\u_div/SumTmp[6][1] ),
	.CO(\u_div/CryTmp[6][2] ),
	.CI(\u_div/CryTmp[6][1] ),
	.B(n17),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_4  (
	.S(\u_div/SumTmp[3][4] ),
	.CO(\u_div/CryTmp[3][5] ),
	.CI(\u_div/CryTmp[3][4] ),
	.B(n14),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(n13),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(n12),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(n11),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_1  (
	.S(\u_div/SumTmp[2][1] ),
	.CO(\u_div/CryTmp[2][2] ),
	.CI(\u_div/CryTmp[2][1] ),
	.B(n17),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_1  (
	.S(\u_div/SumTmp[3][1] ),
	.CO(\u_div/CryTmp[3][2] ),
	.CI(\u_div/CryTmp[3][1] ),
	.B(n17),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_1  (
	.S(\u_div/SumTmp[4][1] ),
	.CO(\u_div/CryTmp[4][2] ),
	.CI(\u_div/CryTmp[4][1] ),
	.B(n17),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_1  (
	.S(\u_div/SumTmp[5][1] ),
	.CO(\u_div/CryTmp[5][2] ),
	.CI(\u_div/CryTmp[5][1] ),
	.B(n17),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(n16),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(n15),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(n14),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_5  (
	.S(\u_div/SumTmp[1][5] ),
	.CO(\u_div/CryTmp[1][6] ),
	.CI(\u_div/CryTmp[1][5] ),
	.B(n13),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_4  (
	.S(\u_div/SumTmp[1][4] ),
	.CO(\u_div/CryTmp[1][5] ),
	.CI(\u_div/CryTmp[1][4] ),
	.B(n14),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_3  (
	.S(\u_div/SumTmp[1][3] ),
	.CO(\u_div/CryTmp[1][4] ),
	.CI(\u_div/CryTmp[1][3] ),
	.B(n15),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_4  (
	.S(\u_div/SumTmp[2][4] ),
	.CO(\u_div/CryTmp[2][5] ),
	.CI(\u_div/CryTmp[2][4] ),
	.B(n14),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_2  (
	.S(\u_div/SumTmp[1][2] ),
	.CO(\u_div/CryTmp[1][3] ),
	.CI(\u_div/CryTmp[1][2] ),
	.B(n16),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_3  (
	.S(\u_div/SumTmp[2][3] ),
	.CO(\u_div/CryTmp[2][4] ),
	.CI(\u_div/CryTmp[2][3] ),
	.B(n15),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_2  (
	.S(\u_div/SumTmp[2][2] ),
	.CO(\u_div/CryTmp[2][3] ),
	.CI(\u_div/CryTmp[2][2] ),
	.B(n16),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_3  (
	.S(\u_div/SumTmp[3][3] ),
	.CO(\u_div/CryTmp[3][4] ),
	.CI(\u_div/CryTmp[3][3] ),
	.B(n15),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_2  (
	.S(\u_div/SumTmp[3][2] ),
	.CO(\u_div/CryTmp[3][3] ),
	.CI(\u_div/CryTmp[3][2] ),
	.B(n16),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_2  (
	.S(\u_div/SumTmp[4][2] ),
	.CO(\u_div/CryTmp[4][3] ),
	.CI(\u_div/CryTmp[4][2] ),
	.B(n16),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(n18),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(\u_div/SumTmp[6][0] ),
	.B(a[6]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(\u_div/SumTmp[5][0] ),
	.B(a[5]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(\u_div/SumTmp[4][0] ),
	.B(a[4]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(\u_div/CryTmp[5][1] ),
	.B(n3),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n3),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n2),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U12 (
	.Y(\u_div/CryTmp[4][1] ),
	.B(n5),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n5),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n4),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U15 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n7),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n6),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n8),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n8),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U20 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(n1),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n1),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U22 (
	.Y(\u_div/SumTmp[1][0] ),
	.B(a[1]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n17),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n16),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n15),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n14),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n13),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n10),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n12),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U30 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(n9),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n9),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(n10),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n11),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U34 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][6] ),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U35 (
	.Y(\u_div/PartRem[2][6] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U36 (
	.Y(\u_div/PartRem[3][5] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U37 (
	.Y(\u_div/PartRem[4][4] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U38 (
	.Y(\u_div/PartRem[5][3] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U39 (
	.Y(\u_div/PartRem[6][2] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][1] ),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U40 (
	.Y(\u_div/PartRem[7][1] ),
	.S0(quotient[7]),
	.B(\u_div/SumTmp[7][0] ),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U41 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][5] ),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U42 (
	.Y(\u_div/PartRem[2][5] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U43 (
	.Y(\u_div/PartRem[3][4] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U44 (
	.Y(\u_div/PartRem[4][3] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][2] ),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U45 (
	.Y(\u_div/PartRem[5][2] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][1] ),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U46 (
	.Y(\u_div/PartRem[6][1] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][0] ),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U47 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][4] ),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U48 (
	.Y(\u_div/PartRem[2][4] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U49 (
	.Y(\u_div/PartRem[3][3] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U50 (
	.Y(\u_div/PartRem[4][2] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][1] ),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U51 (
	.Y(\u_div/PartRem[5][1] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][0] ),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U52 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][3] ),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U53 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U54 (
	.Y(\u_div/PartRem[3][2] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][1] ),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U55 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][0] ),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U56 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][2] ),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U57 (
	.Y(\u_div/PartRem[2][2] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][1] ),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U58 (
	.Y(\u_div/PartRem[3][1] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][0] ),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U59 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][1] ),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U60 (
	.Y(\u_div/PartRem[2][1] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][0] ),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U61 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][0] ),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U62 (
	.Y(quotient[7]),
	.D(n16),
	.C(n17),
	.B(n19),
	.A(\u_div/CryTmp[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U63 (
	.Y(quotient[6]),
	.C(\u_div/CryTmp[6][2] ),
	.B(n16),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U64 (
	.Y(quotient[5]),
	.B(n19),
	.A(\u_div/CryTmp[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U65 (
	.Y(n19),
	.B(n15),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U66 (
	.Y(quotient[4]),
	.B(n20),
	.A(\u_div/CryTmp[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U67 (
	.Y(n20),
	.C(n13),
	.B(n14),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U68 (
	.Y(quotient[3]),
	.C(\u_div/CryTmp[3][5] ),
	.B(n13),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U69 (
	.Y(quotient[2]),
	.B(n21),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(n21),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U71 (
	.Y(quotient[1]),
	.B(n11),
	.A(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n2),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n8),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n3),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n4),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n5),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n6),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n7),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U1 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(n1),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n9),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n7),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n6),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n5),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n4),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n3),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(carry[1]),
	.B(n1),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n8),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n2),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U12 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[0]),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;

   // Module instantiations
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n8),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n9),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n7),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n6),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n5),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n4),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n3),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U10 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(\A1[6] ),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(PRODUCT[1]),
	.B(\ab[0][1] ),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n22),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n21),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n20),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n19),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n18),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n17),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U24 (
	.Y(n11),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U25 (
	.Y(n12),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U26 (
	.Y(n13),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U27 (
	.Y(n14),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n16),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U30 (
	.Y(\SUMB[1][6] ),
	.B(n22),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U31 (
	.Y(\SUMB[1][5] ),
	.B(n21),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(\SUMB[1][4] ),
	.B(n20),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U33 (
	.Y(\SUMB[1][3] ),
	.B(n19),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U34 (
	.Y(\SUMB[1][2] ),
	.B(n18),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][1] ),
	.B(n17),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n31),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n36),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n35),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n34),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n33),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n32),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n38),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n37),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n30),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n24),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n23),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n28),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n29),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n27),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n26),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U51 (
	.Y(n25),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U53 (
	.Y(\ab[7][7] ),
	.B(n23),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U54 (
	.Y(\ab[7][6] ),
	.B(n24),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][5] ),
	.B(n25),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][4] ),
	.B(n26),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][3] ),
	.B(n27),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][2] ),
	.B(n28),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][1] ),
	.B(n29),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][0] ),
	.B(n30),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[6][7] ),
	.B(n32),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[6][6] ),
	.B(n32),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][5] ),
	.B(n32),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][4] ),
	.B(n32),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][3] ),
	.B(n32),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][2] ),
	.B(n32),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][1] ),
	.B(n32),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][0] ),
	.B(n32),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[5][7] ),
	.B(n33),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[5][6] ),
	.B(n33),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][5] ),
	.B(n33),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][4] ),
	.B(n33),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][3] ),
	.B(n33),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][2] ),
	.B(n33),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][1] ),
	.B(n33),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][0] ),
	.B(n33),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[4][7] ),
	.B(n34),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[4][6] ),
	.B(n34),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][5] ),
	.B(n34),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][4] ),
	.B(n34),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][3] ),
	.B(n34),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][2] ),
	.B(n34),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][1] ),
	.B(n34),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][0] ),
	.B(n34),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[3][7] ),
	.B(n35),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[3][6] ),
	.B(n35),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][5] ),
	.B(n35),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][4] ),
	.B(n35),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][3] ),
	.B(n35),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][2] ),
	.B(n35),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][1] ),
	.B(n35),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][0] ),
	.B(n35),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[2][7] ),
	.B(n36),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[2][6] ),
	.B(n36),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][5] ),
	.B(n36),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][4] ),
	.B(n36),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][3] ),
	.B(n36),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][2] ),
	.B(n36),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][1] ),
	.B(n36),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][0] ),
	.B(n36),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[1][7] ),
	.B(n37),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[1][6] ),
	.B(n37),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][5] ),
	.B(n37),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][4] ),
	.B(n37),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][3] ),
	.B(n37),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][2] ),
	.B(n37),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][1] ),
	.B(n37),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][0] ),
	.B(n37),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[0][7] ),
	.B(n38),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[0][6] ),
	.B(n38),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][5] ),
	.B(n38),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][4] ),
	.B(n38),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][3] ),
	.B(n38),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][2] ),
	.B(n38),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][1] ),
	.B(n38),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(PRODUCT[0]),
	.B(n38),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n14,
		n16,
		n13,
		n15,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPERAND_WIDTH8_FUN_WIDTH4_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   // Module instantiations
   AOI21BX2M U2 (
	.Y(n1),
	.B0N(n19),
	.A1(A[12]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n15),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(SUM[7]),
	.B(n8),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n8),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(SUM[6]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n9),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U9 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U10 (
	.Y(SUM[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U11 (
	.Y(SUM[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U12 (
	.Y(SUM[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U13 (
	.Y(SUM[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U14 (
	.Y(SUM[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U15 (
	.Y(SUM[9]),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(SUM[8]),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U18 (
	.Y(n14),
	.B(n17),
	.AN(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(n19),
	.B0(B[12]),
	.A1(n18),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U20 (
	.Y(SUM[12]),
	.C(n18),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U21 (
	.Y(n18),
	.B0N(n22),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U22 (
	.Y(SUM[11]),
	.B(n23),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U23 (
	.Y(n23),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(n20),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U25 (
	.Y(n22),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U26 (
	.Y(n21),
	.B0(n26),
	.A1(n25),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(SUM[10]),
	.B(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U28 (
	.Y(n25),
	.B0(n12),
	.A1N(n13),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U29 (
	.Y(n12),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(n13),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U31 (
	.Y(n10),
	.B0(n17),
	.A1(n16),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n17),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U33 (
	.Y(n16),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U34 (
	.Y(n27),
	.B(n26),
	.AN(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n26),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U36 (
	.Y(n24),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_DIV_MUX (
	IN, 
	OUT, 
	VDD, 
	VSS);
   input [5:0] IN;
   output [7:0] OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n14;
   wire n15;
   wire n16;
   wire n17;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U11 (
	.Y(OUT[1]),
	.C(IN[0]),
	.B(IN[1]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U12 (
	.Y(n6),
	.D(n14),
	.C(n15),
	.B(IN[3]),
	.AN(IN[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U13 (
	.Y(n7),
	.D(n14),
	.C(n15),
	.B(IN[4]),
	.AN(IN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U14 (
	.Y(OUT[2]),
	.C(IN[0]),
	.B(IN[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U15 (
	.Y(OUT[3]),
	.D(IN[4]),
	.C(IN[5]),
	.B(IN[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U16 (
	.Y(n5),
	.C(IN[2]),
	.B(n16),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n15),
	.A(IN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n17),
	.A(IN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n16),
	.A(IN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n14),
	.A(IN[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U21 (
	.Y(OUT[0]),
	.C0(n16),
	.B0(n17),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U22 (
	.Y(n8),
	.D(n15),
	.C(IN[3]),
	.B(IN[4]),
	.A(IN[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(n9),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(OUT[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(OUT[5]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(OUT[6]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(OUT[7]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Clk_Div_WIDTH8_test_0 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN8_SE, 
	UART_SCAN_CLK__L4_N0, 
	UART_SCAN_CLK__L6_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN8_SE;
   input UART_SCAN_CLK__L4_N0;
   input UART_SCAN_CLK__L6_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_div_clk__Exclude_0_NET;
   wire div_clk__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire FE_UNCONNECTED_0;
   wire N0;
   wire div_clk;
   wire flag;
   wire N9;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N19;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n18;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire [7:0] counter;

   assign test_so = flag ;

   // Module instantiations
   DLY3X1M FE_PHC7_div_clk__Exclude_0_NET (
	.Y(FE_PHN7_div_clk__Exclude_0_NET),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M div_clk__Exclude_0 (
	.Y(div_clk__Exclude_0_NET),
	.A(div_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M div_clk_reg (
	.SI(counter[7]),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(div_clk),
	.D(n28),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M flag_reg (
	.SI(FE_PHN7_div_clk__Exclude_0_NET),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(flag),
	.D(n37),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(counter[7]),
	.D(n29),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(n36),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(n34),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(n33),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(n32),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(n31),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(n30),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(n48),
	.SE(FE_OFN8_SE),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(n35),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(n22),
	.B(n21),
	.AN(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U6 (
	.Y(n20),
	.B0(n60),
	.A1N(i_div_ratio[0]),
	.A0(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n60),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U12 (
	.Y(n3),
	.B(i_div_ratio[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U17 (
	.Y(n1),
	.B0N(n3),
	.A1(i_div_ratio[2]),
	.A0(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(N0),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(n23),
	.B(n25),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U20 (
	.Y(n25),
	.B1(flag),
	.B0(N17),
	.A1N(flag),
	.A0(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U21 (
	.Y(n37),
	.B(n24),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(n24),
	.B(n23),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n28),
	.B(n19),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(n19),
	.B(n21),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n29),
	.B1(n22),
	.B0(N31),
	.A1(n21),
	.A0(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n30),
	.B1(n22),
	.B0(N30),
	.A1(n21),
	.A0(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n31),
	.B1(n22),
	.B0(N29),
	.A1(n21),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U28 (
	.Y(n32),
	.B1(n22),
	.B0(N28),
	.A1(n21),
	.A0(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U29 (
	.Y(n33),
	.B1(n22),
	.B0(N27),
	.A1(n21),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U30 (
	.Y(n34),
	.B1(n22),
	.B0(N26),
	.A1(n21),
	.A0(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U31 (
	.Y(n35),
	.B1(n22),
	.B0(N25),
	.A1(n21),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U32 (
	.Y(n36),
	.B1(n22),
	.B0(n48),
	.A1(n21),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U34 (
	.Y(n21),
	.B0(HTIE_LTIEHI_NET),
	.A1N(n27),
	.A0N(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U35 (
	.Y(n27),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U36 (
	.Y(n26),
	.C(i_div_ratio[2]),
	.B(i_div_ratio[3]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n48),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U38 (
	.Y(o_div_clk),
	.S0(N0),
	.B(div_clk),
	.A(UART_SCAN_CLK__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U39 (
	.Y(N9),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U40 (
	.Y(n4),
	.B(i_div_ratio[3]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U41 (
	.Y(N11),
	.B0(n4),
	.A1N(i_div_ratio[3]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U42 (
	.Y(n5),
	.B(LTIE_LTIELO_NET),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U43 (
	.Y(N12),
	.B0(n5),
	.A1N(LTIE_LTIELO_NET),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U44 (
	.Y(n6),
	.B(LTIE_LTIELO_NET),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U45 (
	.Y(N13),
	.B0(n6),
	.A1N(LTIE_LTIELO_NET),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U46 (
	.Y(N14),
	.B(n6),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U47 (
	.Y(N16),
	.C(n6),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U48 (
	.Y(n7),
	.B0(LTIE_LTIELO_NET),
	.A1(n6),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U49 (
	.Y(N15),
	.B(n7),
	.AN(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(n47),
	.B(counter[2]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U51 (
	.Y(n18),
	.B(N9),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U52 (
	.Y(n46),
	.B1(n1),
	.B0(n18),
	.A1(n18),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U53 (
	.Y(n38),
	.B(n48),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U54 (
	.Y(n39),
	.B1(counter[1]),
	.B0(n38),
	.A1(n1),
	.A0(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U55 (
	.Y(n45),
	.C(counter[7]),
	.B(N16),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n43),
	.B(counter[3]),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n42),
	.B(counter[4]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(n41),
	.B(counter[5]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n40),
	.B(counter[6]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U60 (
	.Y(n44),
	.D(n40),
	.C(n41),
	.B(n42),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U61 (
	.Y(N17),
	.D(n44),
	.C(n45),
	.B(n46),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U62 (
	.Y(n49),
	.B(i_div_ratio[1]),
	.AN(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U63 (
	.Y(n53),
	.B1(n49),
	.B0(counter[1]),
	.A1N(i_div_ratio[2]),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U64 (
	.Y(n52),
	.B(counter[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U65 (
	.Y(n50),
	.B(counter[0]),
	.AN(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U66 (
	.Y(n51),
	.B1(n50),
	.B0(i_div_ratio[2]),
	.A1N(counter[1]),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U67 (
	.Y(n59),
	.D(n51),
	.C(n52),
	.B(n53),
	.AN(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U68 (
	.Y(n57),
	.B(counter[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U69 (
	.Y(n56),
	.B(counter[5]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U70 (
	.Y(n55),
	.B(counter[4]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U71 (
	.Y(n54),
	.B(counter[3]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U72 (
	.Y(n58),
	.D(n54),
	.C(n55),
	.B(n56),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(N19),
	.B(n58),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   Clk_Div_WIDTH8_0_DW01_inc_0 add_46 (
	.A({ counter[7],
		counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N31,
		N30,
		N29,
		N28,
		N27,
		N26,
		N25,
		FE_UNCONNECTED_0 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Clk_Div_WIDTH8_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Clk_Div_WIDTH8_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	UART_SCAN_CLK__L4_N0, 
	UART_SCAN_CLK__L6_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input UART_SCAN_CLK__L4_N0;
   input UART_SCAN_CLK__L6_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN6_div_clk__Exclude_0_NET;
   wire div_clk__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire N0;
   wire div_clk;
   wire flag;
   wire N9;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N19;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n18;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire [7:0] counter;

   assign test_so = flag ;

   // Module instantiations
   DLY3X1M FE_PHC6_div_clk__Exclude_0_NET (
	.Y(FE_PHN6_div_clk__Exclude_0_NET),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M div_clk__Exclude_0 (
	.Y(div_clk__Exclude_0_NET),
	.A(div_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M div_clk_reg (
	.SI(counter[7]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(div_clk),
	.D(n70),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M flag_reg (
	.SI(FE_PHN6_div_clk__Exclude_0_NET),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(flag),
	.D(n61),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[7]),
	.D(n69),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(n62),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(n64),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(n65),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(n66),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(n67),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(n68),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(n48),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(n63),
	.CK(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(n76),
	.B(n77),
	.AN(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(N0),
	.A(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U7 (
	.Y(n78),
	.B0(n60),
	.A1N(i_div_ratio[0]),
	.A0(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n60),
	.A(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U17 (
	.Y(n3),
	.B(i_div_ratio[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n75),
	.B(n73),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U19 (
	.Y(n73),
	.B1(flag),
	.B0(N17),
	.A1N(flag),
	.A0(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U20 (
	.Y(n69),
	.B1(n76),
	.B0(N31),
	.A1(n77),
	.A0(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U21 (
	.Y(n68),
	.B1(n76),
	.B0(N30),
	.A1(n77),
	.A0(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U22 (
	.Y(n67),
	.B1(n76),
	.B0(N29),
	.A1(n77),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U23 (
	.Y(n66),
	.B1(n76),
	.B0(N28),
	.A1(n77),
	.A0(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U24 (
	.Y(n65),
	.B1(n76),
	.B0(N27),
	.A1(n77),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n64),
	.B1(n76),
	.B0(N26),
	.A1(n77),
	.A0(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n63),
	.B1(n76),
	.B0(N25),
	.A1(n77),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n62),
	.B1(n76),
	.B0(N24),
	.A1(n77),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U28 (
	.Y(n70),
	.B(n79),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(n79),
	.B(n77),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n61),
	.B(n74),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(n74),
	.B(n75),
	.A(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U32 (
	.Y(n1),
	.B0N(n3),
	.A1(i_div_ratio[2]),
	.A0(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n48),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U35 (
	.Y(n77),
	.B0(HTIE_LTIEHI_NET),
	.A1N(n71),
	.A0N(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U36 (
	.Y(n72),
	.C(i_div_ratio[2]),
	.B(i_div_ratio[3]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U37 (
	.Y(n71),
	.D(i_div_ratio[4]),
	.C(i_div_ratio[5]),
	.B(i_div_ratio[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U38 (
	.Y(o_div_clk),
	.S0(N0),
	.B(div_clk),
	.A(UART_SCAN_CLK__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U39 (
	.Y(N9),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U40 (
	.Y(n4),
	.B(i_div_ratio[3]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U41 (
	.Y(N11),
	.B0(n4),
	.A1N(i_div_ratio[3]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U42 (
	.Y(n5),
	.B(i_div_ratio[4]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U43 (
	.Y(N12),
	.B0(n5),
	.A1N(i_div_ratio[4]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U44 (
	.Y(n6),
	.B(i_div_ratio[5]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U45 (
	.Y(N13),
	.B0(n6),
	.A1N(i_div_ratio[5]),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U46 (
	.Y(N14),
	.B(n6),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U47 (
	.Y(N16),
	.C(n6),
	.B(i_div_ratio[7]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U48 (
	.Y(n7),
	.B0(i_div_ratio[7]),
	.A1(n6),
	.A0(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U49 (
	.Y(N15),
	.B(n7),
	.AN(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(n47),
	.B(counter[2]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U51 (
	.Y(n18),
	.B(N9),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U52 (
	.Y(n46),
	.B1(n1),
	.B0(n18),
	.A1(n18),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U53 (
	.Y(n38),
	.B(n48),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U54 (
	.Y(n39),
	.B1(counter[1]),
	.B0(n38),
	.A1(n1),
	.A0(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U55 (
	.Y(n45),
	.C(counter[7]),
	.B(N16),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n43),
	.B(counter[3]),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n42),
	.B(counter[4]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(n41),
	.B(counter[5]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n40),
	.B(counter[6]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U60 (
	.Y(n44),
	.D(n40),
	.C(n41),
	.B(n42),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U61 (
	.Y(N17),
	.D(n44),
	.C(n45),
	.B(n46),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U62 (
	.Y(n49),
	.B(i_div_ratio[1]),
	.AN(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U63 (
	.Y(n53),
	.B1(n49),
	.B0(counter[1]),
	.A1N(i_div_ratio[2]),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U64 (
	.Y(n52),
	.B(counter[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U65 (
	.Y(n50),
	.B(counter[0]),
	.AN(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U66 (
	.Y(n51),
	.B1(n50),
	.B0(i_div_ratio[2]),
	.A1N(counter[1]),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U67 (
	.Y(n59),
	.D(n51),
	.C(n52),
	.B(n53),
	.AN(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U68 (
	.Y(n57),
	.B(counter[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U69 (
	.Y(n56),
	.B(counter[5]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U70 (
	.Y(n55),
	.B(counter[4]),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U71 (
	.Y(n54),
	.B(counter[3]),
	.A(i_div_ratio[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U72 (
	.Y(n58),
	.D(n54),
	.C(n55),
	.B(n56),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(N19),
	.B(n58),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   Clk_Div_WIDTH8_1_DW01_inc_0 add_46 (
	.A({ counter[7],
		counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N31,
		N30,
		N29,
		N28,
		N27,
		N26,
		N25,
		N24 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Clk_Div_WIDTH8_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 (
	WR_DATA, 
	W_INC, 
	R_INC, 
	W_CLK, 
	W_RST, 
	R_CLK, 
	R_RST, 
	FULL, 
	EMPTY, 
	RD_DATA, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN12_SE, 
	FE_OFN8_SE, 
	FE_OFN9_SE, 
	VDD, 
	VSS);
   input [7:0] WR_DATA;
   input W_INC;
   input R_INC;
   input W_CLK;
   input W_RST;
   input R_CLK;
   input R_RST;
   output FULL;
   output EMPTY;
   output [7:0] RD_DATA;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN12_SE;
   input FE_OFN8_SE;
   input FE_OFN9_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [4:0] WR_PTR;
   wire [4:0] SYNC_WR_PTR;
   wire [4:0] RD_PTR;
   wire [4:0] SYNC_RD_PTR;
   wire [3:0] WR_ADDR;
   wire [3:0] RD_ADDR;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;
   wire SYNOPSYS_UNCONNECTED__3;

   // Module instantiations
   DF_SYNC_ADDRESS_WIDTH4_test_0 DUT0 (
	.CLK(R_CLK),
	.RST(R_RST),
	.ASYNC({ 1'b0,
		WR_PTR[3],
		WR_PTR[2],
		WR_PTR[1],
		WR_PTR[0] }),
	.SYNC({ SYNOPSYS_UNCONNECTED__0,
		SYNC_WR_PTR[3],
		SYNC_WR_PTR[2],
		SYNC_WR_PTR[1],
		SYNC_WR_PTR[0] }),
	.test_si(test_si1),
	.test_se(FE_OFN9_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_ADDRESS_WIDTH4_test_1 DUT1 (
	.CLK(W_CLK),
	.RST(W_RST),
	.ASYNC({ 1'b0,
		RD_PTR[3],
		RD_PTR[2],
		RD_PTR[1],
		RD_PTR[0] }),
	.SYNC({ SYNOPSYS_UNCONNECTED__1,
		SYNC_RD_PTR[3],
		SYNC_RD_PTR[2],
		SYNC_RD_PTR[1],
		SYNC_RD_PTR[0] }),
	.test_si(SYNC_WR_PTR[3]),
	.test_se(FE_OFN9_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_WR_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 DUT2 (
	.W_INC(W_INC),
	.W_CLK(W_CLK),
	.W_RST(W_RST),
	.SYNC_RD_PTR({ 1'b0,
		SYNC_RD_PTR[3],
		SYNC_RD_PTR[2],
		SYNC_RD_PTR[1],
		SYNC_RD_PTR[0] }),
	.WR_ADDR({ WR_ADDR[3],
		WR_ADDR[2],
		WR_ADDR[1],
		WR_ADDR[0] }),
	.WR_PTR({ SYNOPSYS_UNCONNECTED__2,
		WR_PTR[3],
		WR_PTR[2],
		WR_PTR[1],
		WR_PTR[0] }),
	.FULL(FULL),
	.test_se(test_se),
	.FE_OFN9_SE(FE_OFN9_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_RD_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 DUT3 (
	.R_INC(R_INC),
	.R_CLK(R_CLK),
	.R_RST(R_RST),
	.SYNC_WR_PTR({ 1'b0,
		SYNC_WR_PTR[3],
		SYNC_WR_PTR[2],
		SYNC_WR_PTR[1],
		SYNC_WR_PTR[0] }),
	.RD_ADDR({ RD_ADDR[3],
		RD_ADDR[2],
		RD_ADDR[1],
		RD_ADDR[0] }),
	.RD_PTR({ SYNOPSYS_UNCONNECTED__3,
		RD_PTR[3],
		RD_PTR[2],
		RD_PTR[1],
		RD_PTR[0] }),
	.EMPTY(EMPTY),
	.test_si(WR_PTR[3]),
	.test_se(FE_OFN9_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_MEM_CNTRL_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 DUT4 (
	.WR_DATA({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.WR_ADDR({ WR_ADDR[3],
		WR_ADDR[2],
		WR_ADDR[1],
		WR_ADDR[0] }),
	.RD_ADDR({ RD_ADDR[3],
		RD_ADDR[2],
		RD_ADDR[1],
		RD_ADDR[0] }),
	.W_INC(W_INC),
	.R_INC(R_INC),
	.W_CLK(W_CLK),
	.R_CLK(R_CLK),
	.FULL(FULL),
	.RD_DATA({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.test_si2(test_si2),
	.test_si1(RD_PTR[3]),
	.test_so2(test_so2),
	.test_so1(test_so1),
	.test_se(FE_OFN12_SE),
	.FE_OFN8_SE(FE_OFN8_SE),
	.FE_OFN9_SE(FE_OFN9_SE), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_ADDRESS_WIDTH4_test_0 (
	CLK, 
	RST, 
	ASYNC, 
	SYNC, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [4:0] ASYNC;
   output [4:0] SYNC;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [3:0] REG;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[3]  (
	.SI(SYNC[2]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[3]),
	.D(REG[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[2]  (
	.SI(SYNC[1]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[2]),
	.D(REG[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[1]  (
	.SI(SYNC[0]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[1]),
	.D(REG[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[0]  (
	.SI(REG[3]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[0]),
	.D(REG[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3]  (
	.SI(REG[2]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[3]),
	.D(ASYNC[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2]  (
	.SI(REG[1]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[2]),
	.D(ASYNC[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1]  (
	.SI(REG[0]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[1]),
	.D(ASYNC[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(REG[0]),
	.D(ASYNC[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(SYNC[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_ADDRESS_WIDTH4_test_1 (
	CLK, 
	RST, 
	ASYNC, 
	SYNC, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [4:0] ASYNC;
   output [4:0] SYNC;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [3:0] REG;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[2]  (
	.SI(SYNC[1]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[2]),
	.D(REG[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[3]  (
	.SI(SYNC[2]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[3]),
	.D(REG[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[1]  (
	.SI(SYNC[0]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[1]),
	.D(REG[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \SYNC_reg[0]  (
	.SI(REG[3]),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[0]),
	.D(REG[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3]  (
	.SI(REG[2]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[3]),
	.D(ASYNC[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2]  (
	.SI(REG[1]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[2]),
	.D(ASYNC[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1]  (
	.SI(REG[0]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[1]),
	.D(ASYNC[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(REG[0]),
	.D(ASYNC[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(SYNC[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_WR_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 (
	W_INC, 
	W_CLK, 
	W_RST, 
	SYNC_RD_PTR, 
	WR_ADDR, 
	WR_PTR, 
	FULL, 
	test_se, 
	FE_OFN9_SE, 
	VDD, 
	VSS);
   input W_INC;
   input W_CLK;
   input W_RST;
   input [4:0] SYNC_RD_PTR;
   output [3:0] WR_ADDR;
   output [4:0] WR_PTR;
   output FULL;
   input test_se;
   input FE_OFN9_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N110;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n20;
   wire n22;
   wire n24;
   wire n35;
   wire n36;
   wire \add_28/carry[4] ;
   wire \add_28/carry[3] ;
   wire \add_28/carry[2] ;
   wire n4;
   wire n8;
   wire [4:0] WR_PTR_binary;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_reg[2]  (
	.SI(WR_PTR[1]),
	.SE(test_se),
	.RN(W_RST),
	.Q(WR_PTR[2]),
	.D(n22),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_reg[0]  (
	.SI(n36),
	.SE(test_se),
	.RN(W_RST),
	.Q(WR_PTR[0]),
	.D(n35),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_reg[1]  (
	.SI(WR_PTR[0]),
	.SE(test_se),
	.RN(W_RST),
	.Q(WR_PTR[1]),
	.D(n24),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_reg[3]  (
	.SI(WR_PTR[2]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_PTR[3]),
	.D(n20),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_binary_reg[0]  (
	.SI(WR_ADDR[3]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_PTR_binary[0]),
	.D(N34),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_ADDR_reg[3]  (
	.SI(WR_ADDR[2]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_ADDR[3]),
	.D(N33),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_ADDR_reg[2]  (
	.SI(WR_ADDR[1]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_ADDR[2]),
	.D(N32),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_binary_reg[3]  (
	.SI(WR_PTR_binary[2]),
	.SE(test_se),
	.RN(W_RST),
	.Q(N110),
	.D(N37),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_binary_reg[1]  (
	.SI(N25),
	.SE(test_se),
	.RN(W_RST),
	.Q(WR_PTR_binary[1]),
	.D(N35),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_PTR_binary_reg[2]  (
	.SI(WR_PTR_binary[1]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_PTR_binary[2]),
	.D(N36),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_ADDR_reg[0]  (
	.SI(SYNC_RD_PTR[3]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_ADDR[0]),
	.D(N30),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \WR_ADDR_reg[1]  (
	.SI(WR_ADDR[0]),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.Q(WR_ADDR[1]),
	.D(N31),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \WR_PTR_binary_reg[4]  (
	.SI(n8),
	.SE(FE_OFN9_SE),
	.RN(W_RST),
	.QN(n36),
	.Q(WR_PTR_binary[4]),
	.D(N38),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n4),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n9),
	.B(n13),
	.A(W_INC), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U8 (
	.Y(N37),
	.B1(n8),
	.B0(n4),
	.A1N(n4),
	.A0N(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(FULL),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(N32),
	.B(n11),
	.A(WR_ADDR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U11 (
	.Y(n11),
	.B(n12),
	.A(WR_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(N38),
	.B1(n4),
	.B0(n36),
	.A1N(n4),
	.A0N(N29), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U13 (
	.Y(n12),
	.B(n4),
	.A(WR_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U14 (
	.Y(N34),
	.B1(n4),
	.B0(N25),
	.A1(WR_PTR_binary[0]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U15 (
	.Y(N36),
	.B1(n4),
	.B0(N27),
	.A1(WR_PTR_binary[2]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U16 (
	.Y(N35),
	.B1(n4),
	.B0(N26),
	.A1(WR_PTR_binary[1]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(N31),
	.B(n12),
	.A(WR_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(N30),
	.B(n4),
	.A(WR_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(N33),
	.B(n10),
	.A(WR_ADDR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U20 (
	.Y(n10),
	.B(n11),
	.AN(WR_ADDR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U21 (
	.Y(n22),
	.B1(WR_PTR_binary[4]),
	.B0(n5),
	.A1N(WR_PTR[2]),
	.A0N(WR_PTR_binary[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(n5),
	.B(WR_PTR_binary[2]),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U23 (
	.Y(n20),
	.B1(WR_PTR_binary[4]),
	.B0(n8),
	.A1N(WR_PTR[3]),
	.A0N(WR_PTR_binary[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U24 (
	.Y(n24),
	.B1(WR_PTR_binary[4]),
	.B0(n6),
	.A1N(WR_PTR[1]),
	.A0N(WR_PTR_binary[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U25 (
	.Y(n6),
	.B(WR_PTR_binary[2]),
	.A(WR_PTR_binary[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U26 (
	.Y(n35),
	.B1(WR_PTR_binary[4]),
	.B0(n7),
	.A1N(WR_PTR[0]),
	.A0N(WR_PTR_binary[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U27 (
	.Y(n7),
	.B(WR_PTR_binary[1]),
	.A(WR_PTR_binary[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n8),
	.A(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U29 (
	.S(N27),
	.CO(\add_28/carry[3] ),
	.B(\add_28/carry[2] ),
	.A(WR_PTR_binary[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U30 (
	.S(N26),
	.CO(\add_28/carry[2] ),
	.B(WR_PTR_binary[0]),
	.A(WR_PTR_binary[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U31 (
	.S(N28),
	.CO(\add_28/carry[4] ),
	.B(\add_28/carry[3] ),
	.A(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U32 (
	.Y(n13),
	.D(n16),
	.C(n15),
	.B(n14),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n14),
	.B(SYNC_RD_PTR[3]),
	.A(WR_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(n16),
	.B(n18),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U49 (
	.Y(n15),
	.B(SYNC_RD_PTR[2]),
	.A(WR_PTR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n17),
	.B(SYNC_RD_PTR[0]),
	.A(WR_PTR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n18),
	.B(SYNC_RD_PTR[1]),
	.A(WR_PTR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U52 (
	.Y(N25),
	.A(WR_PTR_binary[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(N29),
	.B(WR_PTR_binary[4]),
	.A(\add_28/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(WR_PTR[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_RD_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 (
	R_INC, 
	R_CLK, 
	R_RST, 
	SYNC_WR_PTR, 
	RD_ADDR, 
	RD_PTR, 
	EMPTY, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input R_INC;
   input R_CLK;
   input R_RST;
   input [4:0] SYNC_WR_PTR;
   output [3:0] RD_ADDR;
   output [4:0] RD_PTR;
   output EMPTY;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N110;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n18;
   wire n20;
   wire n22;
   wire n29;
   wire n30;
   wire n31;
   wire \add_28/carry[4] ;
   wire \add_28/carry[3] ;
   wire \add_28/carry[2] ;
   wire n8;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire [4:0] RD_PTR_binary;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_ADDR_reg[3]  (
	.SI(n31),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_ADDR[3]),
	.D(N33),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_binary_reg[0]  (
	.SI(RD_ADDR[3]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR_binary[0]),
	.D(N34),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_ADDR_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_ADDR[0]),
	.D(N30),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_binary_reg[3]  (
	.SI(RD_PTR_binary[2]),
	.SE(test_se),
	.RN(R_RST),
	.Q(N110),
	.D(N37),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_binary_reg[1]  (
	.SI(N25),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR_binary[1]),
	.D(N35),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_binary_reg[2]  (
	.SI(RD_PTR_binary[1]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR_binary[2]),
	.D(N36),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_ADDR_reg[1]  (
	.SI(RD_ADDR[0]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_ADDR[1]),
	.D(N31),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_reg[2]  (
	.SI(RD_PTR[1]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR[2]),
	.D(n20),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_reg[3]  (
	.SI(RD_PTR[2]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR[3]),
	.D(n18),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_reg[0]  (
	.SI(n30),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR[0]),
	.D(n29),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RD_PTR_reg[1]  (
	.SI(RD_PTR[0]),
	.SE(test_se),
	.RN(R_RST),
	.Q(RD_PTR[1]),
	.D(n22),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \RD_PTR_binary_reg[4]  (
	.SI(n37),
	.SE(test_se),
	.RN(R_RST),
	.QN(n30),
	.Q(RD_PTR_binary[4]),
	.D(N38),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \RD_ADDR_reg[2]  (
	.SI(RD_ADDR[1]),
	.SE(test_se),
	.RN(R_RST),
	.QN(n31),
	.Q(RD_ADDR[2]),
	.D(N32),
	.CK(R_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U7 (
	.Y(N37),
	.B1(n37),
	.B0(n36),
	.A1N(n36),
	.A0N(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n36),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n11),
	.B(n12),
	.A(RD_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U10 (
	.Y(n9),
	.B(R_INC),
	.AN(EMPTY), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U11 (
	.Y(N38),
	.B1(n36),
	.B0(n30),
	.A1N(n36),
	.A0N(N29), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U12 (
	.Y(n12),
	.B(n36),
	.A(RD_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U13 (
	.Y(N34),
	.B1(n36),
	.B0(N25),
	.A1(RD_PTR_binary[0]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U14 (
	.Y(N36),
	.B1(n36),
	.B0(N27),
	.A1(RD_PTR_binary[2]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U15 (
	.Y(N35),
	.B1(n36),
	.B0(N26),
	.A1(RD_PTR_binary[1]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(N31),
	.B(n12),
	.A(RD_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(N33),
	.B(n10),
	.A(RD_ADDR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(n10),
	.B(n11),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(N30),
	.B(n36),
	.A(RD_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U20 (
	.Y(N32),
	.B(n31),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U21 (
	.Y(n20),
	.B1(RD_PTR_binary[4]),
	.B0(n5),
	.A1N(RD_PTR_binary[4]),
	.A0N(RD_PTR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(n5),
	.B(RD_PTR_binary[2]),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U23 (
	.Y(n18),
	.B1(RD_PTR_binary[4]),
	.B0(n37),
	.A1N(RD_PTR_binary[4]),
	.A0N(RD_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U24 (
	.Y(n22),
	.B1(RD_PTR_binary[4]),
	.B0(n6),
	.A1N(RD_PTR_binary[4]),
	.A0N(RD_PTR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U25 (
	.Y(n6),
	.B(RD_PTR_binary[2]),
	.A(RD_PTR_binary[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U26 (
	.Y(n29),
	.B1(RD_PTR_binary[4]),
	.B0(n7),
	.A1N(RD_PTR_binary[4]),
	.A0N(RD_PTR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U41 (
	.Y(n7),
	.B(RD_PTR_binary[1]),
	.A(RD_PTR_binary[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n37),
	.A(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U43 (
	.S(N27),
	.CO(\add_28/carry[3] ),
	.B(\add_28/carry[2] ),
	.A(RD_PTR_binary[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U44 (
	.S(N26),
	.CO(\add_28/carry[2] ),
	.B(RD_PTR_binary[0]),
	.A(RD_PTR_binary[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U45 (
	.S(N28),
	.CO(\add_28/carry[4] ),
	.B(\add_28/carry[3] ),
	.A(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U46 (
	.Y(N25),
	.A(RD_PTR_binary[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(N29),
	.B(RD_PTR_binary[4]),
	.A(\add_28/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U48 (
	.Y(n32),
	.B(RD_PTR[2]),
	.A(SYNC_WR_PTR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U49 (
	.Y(n8),
	.B(RD_PTR[3]),
	.A(SYNC_WR_PTR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U50 (
	.Y(n35),
	.B(n8),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n34),
	.B(RD_PTR[1]),
	.A(SYNC_WR_PTR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n33),
	.B(RD_PTR[0]),
	.A(SYNC_WR_PTR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U53 (
	.Y(EMPTY),
	.D(n33),
	.C(LTIE_LTIELO_NET),
	.B(n34),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(RD_PTR[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_MEM_CNTRL_DATA_WIDTH8_ADDRESS_WIDTH4_test_1 (
	WR_DATA, 
	WR_ADDR, 
	RD_ADDR, 
	W_INC, 
	R_INC, 
	W_CLK, 
	R_CLK, 
	FULL, 
	RD_DATA, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN8_SE, 
	FE_OFN9_SE, 
	VDD, 
	VSS);
   input [7:0] WR_DATA;
   input [3:0] WR_ADDR;
   input [3:0] RD_ADDR;
   input W_INC;
   input R_INC;
   input W_CLK;
   input R_CLK;
   input FULL;
   output [7:0] RD_DATA;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN8_SE;
   input FE_OFN9_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N9;
   wire N10;
   wire N11;
   wire \MEM[7][7] ;
   wire \MEM[7][6] ;
   wire \MEM[7][5] ;
   wire \MEM[7][4] ;
   wire \MEM[7][3] ;
   wire \MEM[7][2] ;
   wire \MEM[7][1] ;
   wire \MEM[7][0] ;
   wire \MEM[6][7] ;
   wire \MEM[6][6] ;
   wire \MEM[6][5] ;
   wire \MEM[6][4] ;
   wire \MEM[6][3] ;
   wire \MEM[6][2] ;
   wire \MEM[6][1] ;
   wire \MEM[6][0] ;
   wire \MEM[5][7] ;
   wire \MEM[5][6] ;
   wire \MEM[5][5] ;
   wire \MEM[5][4] ;
   wire \MEM[5][3] ;
   wire \MEM[5][2] ;
   wire \MEM[5][1] ;
   wire \MEM[5][0] ;
   wire \MEM[4][7] ;
   wire \MEM[4][6] ;
   wire \MEM[4][5] ;
   wire \MEM[4][4] ;
   wire \MEM[4][3] ;
   wire \MEM[4][2] ;
   wire \MEM[4][1] ;
   wire \MEM[4][0] ;
   wire \MEM[3][7] ;
   wire \MEM[3][6] ;
   wire \MEM[3][5] ;
   wire \MEM[3][4] ;
   wire \MEM[3][3] ;
   wire \MEM[3][2] ;
   wire \MEM[3][1] ;
   wire \MEM[3][0] ;
   wire \MEM[2][7] ;
   wire \MEM[2][6] ;
   wire \MEM[2][5] ;
   wire \MEM[2][4] ;
   wire \MEM[2][3] ;
   wire \MEM[2][2] ;
   wire \MEM[2][1] ;
   wire \MEM[2][0] ;
   wire \MEM[1][7] ;
   wire \MEM[1][6] ;
   wire \MEM[1][5] ;
   wire \MEM[1][4] ;
   wire \MEM[1][3] ;
   wire \MEM[1][2] ;
   wire \MEM[1][1] ;
   wire \MEM[1][0] ;
   wire \MEM[0][7] ;
   wire \MEM[0][6] ;
   wire \MEM[0][5] ;
   wire \MEM[0][4] ;
   wire \MEM[0][3] ;
   wire \MEM[0][2] ;
   wire \MEM[0][1] ;
   wire \MEM[0][0] ;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;

   assign N9 = RD_ADDR[0] ;
   assign N10 = RD_ADDR[1] ;
   assign N11 = RD_ADDR[2] ;
   assign test_so2 = \MEM[7][7]  ;
   assign test_so1 = \MEM[0][3]  ;

   // Module instantiations
   SDFFQX2M \MEM_reg[5][6]  (
	.SI(\MEM[5][5] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[5][6] ),
	.D(n133),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[5][5]  (
	.SI(\MEM[5][4] ),
	.SE(test_se),
	.Q(\MEM[5][5] ),
	.D(n132),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[5][4]  (
	.SI(\MEM[5][3] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[5][4] ),
	.D(n131),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[5][3]  (
	.SI(\MEM[5][2] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[5][3] ),
	.D(n130),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[5][2]  (
	.SI(\MEM[5][1] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[5][2] ),
	.D(n129),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[5][1]  (
	.SI(\MEM[5][0] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[5][1] ),
	.D(n128),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[5][0]  (
	.SI(\MEM[4][7] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[5][0] ),
	.D(n127),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][7]  (
	.SI(\MEM[1][6] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][7] ),
	.D(n102),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][6]  (
	.SI(\MEM[1][5] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][6] ),
	.D(n101),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][5]  (
	.SI(\MEM[1][4] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][5] ),
	.D(n100),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][4]  (
	.SI(\MEM[1][3] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][4] ),
	.D(n99),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][3]  (
	.SI(\MEM[1][2] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][3] ),
	.D(n98),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][2]  (
	.SI(\MEM[1][1] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][2] ),
	.D(n97),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][1]  (
	.SI(\MEM[1][0] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][1] ),
	.D(n96),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[1][0]  (
	.SI(\MEM[0][7] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[1][0] ),
	.D(n95),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][7]  (
	.SI(\MEM[7][6] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][7] ),
	.D(n150),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][6]  (
	.SI(\MEM[7][5] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][6] ),
	.D(n149),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][5]  (
	.SI(\MEM[7][4] ),
	.SE(test_se),
	.Q(\MEM[7][5] ),
	.D(n148),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][4]  (
	.SI(\MEM[7][3] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][4] ),
	.D(n147),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][3]  (
	.SI(\MEM[7][2] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][3] ),
	.D(n146),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][2]  (
	.SI(\MEM[7][1] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][2] ),
	.D(n145),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][1]  (
	.SI(\MEM[7][0] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][1] ),
	.D(n144),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[7][0]  (
	.SI(\MEM[6][7] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[7][0] ),
	.D(n143),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][7]  (
	.SI(\MEM[3][6] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][7] ),
	.D(n118),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][6]  (
	.SI(\MEM[3][5] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][6] ),
	.D(n117),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][5]  (
	.SI(\MEM[3][4] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][5] ),
	.D(n116),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][4]  (
	.SI(\MEM[3][3] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][4] ),
	.D(n115),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][3]  (
	.SI(\MEM[3][2] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][3] ),
	.D(n114),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][2]  (
	.SI(\MEM[3][1] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][2] ),
	.D(n113),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][1]  (
	.SI(\MEM[3][0] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][1] ),
	.D(n112),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[3][0]  (
	.SI(\MEM[2][7] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[3][0] ),
	.D(n111),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][7]  (
	.SI(\MEM[6][6] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[6][7] ),
	.D(n142),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][6]  (
	.SI(\MEM[6][5] ),
	.SE(test_se),
	.Q(\MEM[6][6] ),
	.D(n141),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][5]  (
	.SI(\MEM[6][4] ),
	.SE(test_se),
	.Q(\MEM[6][5] ),
	.D(n140),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][4]  (
	.SI(\MEM[6][3] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[6][4] ),
	.D(n139),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][3]  (
	.SI(\MEM[6][2] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[6][3] ),
	.D(n138),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][2]  (
	.SI(\MEM[6][1] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[6][2] ),
	.D(n137),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][1]  (
	.SI(\MEM[6][0] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[6][1] ),
	.D(n136),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[6][0]  (
	.SI(\MEM[5][7] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[6][0] ),
	.D(n135),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][7]  (
	.SI(\MEM[2][6] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][7] ),
	.D(n110),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][6]  (
	.SI(\MEM[2][5] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][6] ),
	.D(n109),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][5]  (
	.SI(\MEM[2][4] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][5] ),
	.D(n108),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][4]  (
	.SI(\MEM[2][3] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][4] ),
	.D(n107),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][3]  (
	.SI(\MEM[2][2] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][3] ),
	.D(n106),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][2]  (
	.SI(\MEM[2][1] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][2] ),
	.D(n105),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][1]  (
	.SI(\MEM[2][0] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][1] ),
	.D(n104),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[2][0]  (
	.SI(\MEM[1][7] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[2][0] ),
	.D(n103),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][7]  (
	.SI(\MEM[4][6] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][7] ),
	.D(n126),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][6]  (
	.SI(\MEM[4][5] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][6] ),
	.D(n125),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][5]  (
	.SI(\MEM[4][4] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][5] ),
	.D(n124),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][4]  (
	.SI(\MEM[4][3] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][4] ),
	.D(n123),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][3]  (
	.SI(\MEM[4][2] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][3] ),
	.D(n122),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][2]  (
	.SI(\MEM[4][1] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][2] ),
	.D(n121),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][1]  (
	.SI(\MEM[4][0] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[4][1] ),
	.D(n120),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[4][0]  (
	.SI(\MEM[3][7] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[4][0] ),
	.D(n119),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][7]  (
	.SI(\MEM[0][6] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][7] ),
	.D(n94),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][6]  (
	.SI(\MEM[0][5] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][6] ),
	.D(n93),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][5]  (
	.SI(\MEM[0][4] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][5] ),
	.D(n92),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][4]  (
	.SI(test_si2),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][4] ),
	.D(n91),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][3]  (
	.SI(\MEM[0][2] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][3] ),
	.D(n90),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][2]  (
	.SI(\MEM[0][1] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][2] ),
	.D(n89),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][1]  (
	.SI(\MEM[0][0] ),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][1] ),
	.D(n88),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \MEM_reg[0][0]  (
	.SI(test_si1),
	.SE(FE_OFN9_SE),
	.Q(\MEM[0][0] ),
	.D(n87),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX1M \MEM_reg[5][7]  (
	.SI(\MEM[5][6] ),
	.SE(FE_OFN8_SE),
	.Q(\MEM[5][7] ),
	.D(n134),
	.CK(W_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U67 (
	.Y(n76),
	.B(WR_ADDR[2]),
	.AN(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U71 (
	.Y(n81),
	.C(n82),
	.B(n172),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U72 (
	.Y(n75),
	.C(n76),
	.B(n172),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U73 (
	.Y(n78),
	.C(WR_ADDR[1]),
	.B(n171),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U74 (
	.Y(n79),
	.C(WR_ADDR[1]),
	.B(n76),
	.A(WR_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U75 (
	.Y(n77),
	.C(WR_ADDR[0]),
	.B(n172),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U76 (
	.Y(n163),
	.A(WR_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U77 (
	.Y(n164),
	.A(WR_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U78 (
	.Y(n165),
	.A(WR_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(n166),
	.A(WR_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U80 (
	.Y(n167),
	.A(WR_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U81 (
	.Y(n168),
	.A(WR_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U82 (
	.Y(n169),
	.A(WR_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U83 (
	.Y(n170),
	.A(WR_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n87),
	.B1(n163),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n88),
	.B1(n164),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n89),
	.B1(n165),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n90),
	.B1(n166),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n91),
	.B1(n167),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n92),
	.B1(n168),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n93),
	.B1(n169),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n94),
	.B1(n170),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U92 (
	.Y(n103),
	.B1(n78),
	.B0(n163),
	.A1N(n78),
	.A0N(\MEM[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U93 (
	.Y(n104),
	.B1(n78),
	.B0(n164),
	.A1N(n78),
	.A0N(\MEM[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U94 (
	.Y(n105),
	.B1(n78),
	.B0(n165),
	.A1N(n78),
	.A0N(\MEM[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n106),
	.B1(n78),
	.B0(n166),
	.A1N(n78),
	.A0N(\MEM[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U96 (
	.Y(n107),
	.B1(n78),
	.B0(n167),
	.A1N(n78),
	.A0N(\MEM[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U97 (
	.Y(n108),
	.B1(n78),
	.B0(n168),
	.A1N(n78),
	.A0N(\MEM[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U98 (
	.Y(n109),
	.B1(n78),
	.B0(n169),
	.A1N(n78),
	.A0N(\MEM[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U99 (
	.Y(n110),
	.B1(n78),
	.B0(n170),
	.A1N(n78),
	.A0N(\MEM[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n111),
	.B1(n79),
	.B0(n163),
	.A1N(n79),
	.A0N(\MEM[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n112),
	.B1(n79),
	.B0(n164),
	.A1N(n79),
	.A0N(\MEM[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n113),
	.B1(n79),
	.B0(n165),
	.A1N(n79),
	.A0N(\MEM[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n114),
	.B1(n79),
	.B0(n166),
	.A1N(n79),
	.A0N(\MEM[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n115),
	.B1(n79),
	.B0(n167),
	.A1N(n79),
	.A0N(\MEM[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U105 (
	.Y(n116),
	.B1(n79),
	.B0(n168),
	.A1N(n79),
	.A0N(\MEM[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U106 (
	.Y(n117),
	.B1(n79),
	.B0(n169),
	.A1N(n79),
	.A0N(\MEM[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U107 (
	.Y(n118),
	.B1(n79),
	.B0(n170),
	.A1N(n79),
	.A0N(\MEM[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U108 (
	.Y(n95),
	.B1(n77),
	.B0(n163),
	.A1N(n77),
	.A0N(\MEM[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U109 (
	.Y(n96),
	.B1(n77),
	.B0(n164),
	.A1N(n77),
	.A0N(\MEM[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U110 (
	.Y(n97),
	.B1(n77),
	.B0(n165),
	.A1N(n77),
	.A0N(\MEM[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U111 (
	.Y(n98),
	.B1(n77),
	.B0(n166),
	.A1N(n77),
	.A0N(\MEM[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U112 (
	.Y(n99),
	.B1(n77),
	.B0(n167),
	.A1N(n77),
	.A0N(\MEM[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U113 (
	.Y(n100),
	.B1(n77),
	.B0(n168),
	.A1N(n77),
	.A0N(\MEM[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U114 (
	.Y(n101),
	.B1(n77),
	.B0(n169),
	.A1N(n77),
	.A0N(\MEM[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U115 (
	.Y(n102),
	.B1(n77),
	.B0(n170),
	.A1N(n77),
	.A0N(\MEM[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U116 (
	.Y(n119),
	.B1(n81),
	.B0(n163),
	.A1N(n81),
	.A0N(\MEM[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U117 (
	.Y(n120),
	.B1(n81),
	.B0(n164),
	.A1N(n81),
	.A0N(\MEM[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n121),
	.B1(n81),
	.B0(n165),
	.A1N(n81),
	.A0N(\MEM[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n122),
	.B1(n81),
	.B0(n166),
	.A1N(n81),
	.A0N(\MEM[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n123),
	.B1(n81),
	.B0(n167),
	.A1N(n81),
	.A0N(\MEM[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n124),
	.B1(n81),
	.B0(n168),
	.A1N(n81),
	.A0N(\MEM[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n125),
	.B1(n81),
	.B0(n169),
	.A1N(n81),
	.A0N(\MEM[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n126),
	.B1(n81),
	.B0(n170),
	.A1N(n81),
	.A0N(\MEM[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n127),
	.B1(n83),
	.B0(n163),
	.A1N(n83),
	.A0N(\MEM[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U125 (
	.Y(n128),
	.B1(n83),
	.B0(n164),
	.A1N(n83),
	.A0N(\MEM[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U126 (
	.Y(n129),
	.B1(n83),
	.B0(n165),
	.A1N(n83),
	.A0N(\MEM[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U127 (
	.Y(n130),
	.B1(n83),
	.B0(n166),
	.A1N(n83),
	.A0N(\MEM[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U128 (
	.Y(n131),
	.B1(n83),
	.B0(n167),
	.A1N(n83),
	.A0N(\MEM[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U129 (
	.Y(n132),
	.B1(n83),
	.B0(n168),
	.A1N(n83),
	.A0N(\MEM[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U130 (
	.Y(n133),
	.B1(n83),
	.B0(n169),
	.A1N(n83),
	.A0N(\MEM[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U131 (
	.Y(n134),
	.B1(n83),
	.B0(n170),
	.A1N(n83),
	.A0N(\MEM[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U132 (
	.Y(n135),
	.B1(n84),
	.B0(n163),
	.A1N(n84),
	.A0N(\MEM[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U133 (
	.Y(n136),
	.B1(n84),
	.B0(n164),
	.A1N(n84),
	.A0N(\MEM[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U134 (
	.Y(n137),
	.B1(n84),
	.B0(n165),
	.A1N(n84),
	.A0N(\MEM[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U135 (
	.Y(n138),
	.B1(n84),
	.B0(n166),
	.A1N(n84),
	.A0N(\MEM[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n139),
	.B1(n84),
	.B0(n167),
	.A1N(n84),
	.A0N(\MEM[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n140),
	.B1(n84),
	.B0(n168),
	.A1N(n84),
	.A0N(\MEM[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n141),
	.B1(n84),
	.B0(n169),
	.A1N(n84),
	.A0N(\MEM[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n142),
	.B1(n84),
	.B0(n170),
	.A1N(n84),
	.A0N(\MEM[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n143),
	.B1(n85),
	.B0(n163),
	.A1N(n85),
	.A0N(\MEM[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n144),
	.B1(n85),
	.B0(n164),
	.A1N(n85),
	.A0N(\MEM[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n145),
	.B1(n85),
	.B0(n165),
	.A1N(n85),
	.A0N(\MEM[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n146),
	.B1(n85),
	.B0(n166),
	.A1N(n85),
	.A0N(\MEM[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n147),
	.B1(n85),
	.B0(n167),
	.A1N(n85),
	.A0N(\MEM[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n148),
	.B1(n85),
	.B0(n168),
	.A1N(n85),
	.A0N(\MEM[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n149),
	.B1(n85),
	.B0(n169),
	.A1N(n85),
	.A0N(\MEM[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n150),
	.B1(n85),
	.B0(n170),
	.A1N(n85),
	.A0N(\MEM[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U148 (
	.Y(n82),
	.B(n80),
	.A(WR_ADDR[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U149 (
	.Y(n83),
	.C(n82),
	.B(n172),
	.A(WR_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U150 (
	.Y(n84),
	.C(n82),
	.B(n171),
	.A(WR_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U151 (
	.Y(n85),
	.C(n82),
	.B(WR_ADDR[0]),
	.A(WR_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U152 (
	.Y(n80),
	.B(W_INC),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U153 (
	.Y(n86),
	.B(FULL),
	.A(WR_ADDR[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U154 (
	.Y(n172),
	.A(WR_ADDR[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U155 (
	.Y(n171),
	.A(WR_ADDR[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U156 (
	.Y(RD_DATA[0]),
	.S0(N11),
	.B(n66),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U157 (
	.Y(n67),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][0] ),
	.C(\MEM[2][0] ),
	.B(\MEM[1][0] ),
	.A(\MEM[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U158 (
	.Y(n66),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][0] ),
	.C(\MEM[6][0] ),
	.B(\MEM[5][0] ),
	.A(\MEM[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U159 (
	.Y(RD_DATA[4]),
	.S0(N11),
	.B(n74),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U160 (
	.Y(n151),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][4] ),
	.C(\MEM[2][4] ),
	.B(\MEM[1][4] ),
	.A(\MEM[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U161 (
	.Y(n74),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][4] ),
	.C(\MEM[6][4] ),
	.B(\MEM[5][4] ),
	.A(\MEM[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U162 (
	.Y(RD_DATA[1]),
	.S0(N11),
	.B(n68),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U163 (
	.Y(n69),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][1] ),
	.C(\MEM[2][1] ),
	.B(\MEM[1][1] ),
	.A(\MEM[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U164 (
	.Y(n68),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][1] ),
	.C(\MEM[6][1] ),
	.B(\MEM[5][1] ),
	.A(\MEM[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U165 (
	.Y(RD_DATA[2]),
	.S0(N11),
	.B(n70),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U166 (
	.Y(n71),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][2] ),
	.C(\MEM[2][2] ),
	.B(\MEM[1][2] ),
	.A(\MEM[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U167 (
	.Y(n70),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][2] ),
	.C(\MEM[6][2] ),
	.B(\MEM[5][2] ),
	.A(\MEM[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U168 (
	.Y(RD_DATA[3]),
	.S0(N11),
	.B(n72),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U169 (
	.Y(n73),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][3] ),
	.C(\MEM[2][3] ),
	.B(\MEM[1][3] ),
	.A(\MEM[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U170 (
	.Y(n72),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][3] ),
	.C(\MEM[6][3] ),
	.B(\MEM[5][3] ),
	.A(\MEM[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U171 (
	.Y(RD_DATA[5]),
	.S0(N11),
	.B(n152),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U172 (
	.Y(n153),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][5] ),
	.C(\MEM[2][5] ),
	.B(\MEM[1][5] ),
	.A(\MEM[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U173 (
	.Y(n152),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][5] ),
	.C(\MEM[6][5] ),
	.B(\MEM[5][5] ),
	.A(\MEM[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U174 (
	.Y(RD_DATA[6]),
	.S0(N11),
	.B(n154),
	.A(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U175 (
	.Y(n155),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][6] ),
	.C(\MEM[2][6] ),
	.B(\MEM[1][6] ),
	.A(\MEM[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U176 (
	.Y(n154),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][6] ),
	.C(\MEM[6][6] ),
	.B(\MEM[5][6] ),
	.A(\MEM[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U177 (
	.Y(RD_DATA[7]),
	.S0(N11),
	.B(n156),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U178 (
	.Y(n157),
	.S1(N10),
	.S0(n159),
	.D(\MEM[3][7] ),
	.C(\MEM[2][7] ),
	.B(\MEM[1][7] ),
	.A(\MEM[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U179 (
	.Y(n156),
	.S1(N10),
	.S0(n158),
	.D(\MEM[7][7] ),
	.C(\MEM[6][7] ),
	.B(\MEM[5][7] ),
	.A(\MEM[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U180 (
	.Y(n158),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U181 (
	.Y(n159),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GEN_test_1 (
	CLK, 
	RST, 
	LVL_SIG, 
	PULSE_SIG, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN9_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input LVL_SIG;
   output PULSE_SIG;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN9_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FLOP_OUT;
   wire FLOP_IN;

   assign test_so = FLOP_OUT ;

   // Module instantiations
   SDFFRQX2M FLOP_IN_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(FLOP_IN),
	.D(LVL_SIG),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M FLOP_OUT_reg (
	.SI(FLOP_IN),
	.SE(FE_OFN9_SE),
	.RN(RST),
	.Q(FLOP_OUT),
	.D(FLOP_IN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(PULSE_SIG),
	.B(FLOP_OUT),
	.AN(FLOP_IN), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_RX_test_1 (
	clk, 
	rst, 
	rx_in, 
	par_en, 
	par_typ, 
	prescale, 
	data_valid, 
	par_error, 
	stp_error, 
	p_data, 
	test_si, 
	test_se, 
	FE_OFN3_SYNC_UART_SCAN_RST, 
	FE_OFN12_SE, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input rx_in;
   input par_en;
   input par_typ;
   input [5:0] prescale;
   output data_valid;
   output par_error;
   output stp_error;
   output [7:0] p_data;
   input test_si;
   input test_se;
   input FE_OFN3_SYNC_UART_SCAN_RST;
   input FE_OFN12_SE;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PT1_;
   wire FE_UNCONNECTED_0;
   wire str_glitch;
   wire par_chk_en;
   wire str_chk_en;
   wire stp_chk_en;
   wire counter_en;
   wire deser_en;
   wire sampled_bit;
   wire n3;
   wire n4;
   wire [3:0] bit_count;
   wire [4:0] edge_count;

   // Module instantiations
   fsm_test_1 DUT0 (
	.clk(clk),
	.rst(rst),
	.rx_in(rx_in),
	.par_en(par_en),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.par_error(par_error),
	.str_glitch(str_glitch),
	.stp_error(stp_error),
	.prescale({ prescale[5],
		prescale[4],
		prescale[3],
		prescale[2],
		prescale[1],
		prescale[0] }),
	.par_chk_en(par_chk_en),
	.str_chk_en(str_chk_en),
	.stp_chk_en(stp_chk_en),
	.data_sample_en(FE_PT1_),
	.counter_en(counter_en),
	.deser_en(deser_en),
	.data_valid(data_valid),
	.test_si(test_si),
	.test_so(n4),
	.test_se(FE_OFN12_SE),
	.FE_OFN3_SYNC_UART_SCAN_RST(FE_OFN3_SYNC_UART_SCAN_RST),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   counter_test_1 DUT1 (
	.clk(clk),
	.rst(rst),
	.counter_en(counter_en),
	.prescale({ prescale[5],
		prescale[4],
		prescale[3],
		prescale[2],
		prescale[1],
		prescale[0] }),
	.par_en(par_en),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.test_si(n4),
	.test_se(FE_OFN12_SE),
	.FE_OFN3_SYNC_UART_SCAN_RST(FE_OFN3_SYNC_UART_SCAN_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   data_sampling_test_1 DUT2 (
	.clk(clk),
	.rst(rst),
	.rx_in(rx_in),
	.prescale({ prescale[5],
		prescale[4],
		prescale[3],
		prescale[2],
		prescale[1],
		prescale[0] }),
	.edge_count({ edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.data_sample_en(counter_en),
	.sampled_bit(sampled_bit),
	.test_so(n3),
	.test_se(FE_OFN12_SE),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_check_test_1 DUT3 (
	.clk(clk),
	.rst(rst),
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.par_typ(par_typ),
	.par_chk_en(par_chk_en),
	.sampled_bit(sampled_bit),
	.par_error(par_error),
	.test_si(n3),
	.test_se(FE_OFN12_SE),
	.FE_OFN3_SYNC_UART_SCAN_RST(FE_OFN3_SYNC_UART_SCAN_RST),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   start_check_test_1 DUT4 (
	.clk(clk),
	.rst(FE_OFN3_SYNC_UART_SCAN_RST),
	.str_chk_en(str_chk_en),
	.sampled_bit(sampled_bit),
	.str_glitch(str_glitch),
	.test_si(par_error),
	.test_se(FE_OFN12_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   stop_check_test_1 DUT5 (
	.clk(clk),
	.rst(FE_OFN3_SYNC_UART_SCAN_RST),
	.stp_chk_en(stp_chk_en),
	.sampled_bit(sampled_bit),
	.stp_error(stp_error),
	.test_si(str_glitch),
	.test_se(FE_OFN12_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_test_1 DUT6 (
	.clk(clk),
	.rst(rst),
	.deser_en(deser_en),
	.sampled_bit(sampled_bit),
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.test_si(stp_error),
	.test_se(test_se),
	.FE_OFN3_SYNC_UART_SCAN_RST(FE_OFN3_SYNC_UART_SCAN_RST),
	.FE_OFN12_SE(FE_OFN12_SE),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module fsm_test_1 (
	clk, 
	rst, 
	rx_in, 
	par_en, 
	bit_count, 
	edge_count, 
	par_error, 
	str_glitch, 
	stp_error, 
	prescale, 
	par_chk_en, 
	str_chk_en, 
	stp_chk_en, 
	data_sample_en, 
	counter_en, 
	deser_en, 
	data_valid, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN3_SYNC_UART_SCAN_RST, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input rx_in;
   input par_en;
   input [3:0] bit_count;
   input [4:0] edge_count;
   input par_error;
   input str_glitch;
   input stp_error;
   input [5:0] prescale;
   output par_chk_en;
   output str_chk_en;
   output stp_chk_en;
   output data_sample_en;
   output counter_en;
   output deser_en;
   output data_valid;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN3_SYNC_UART_SCAN_RST;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n30;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire \r91/EQ ;
   wire \r91/B[0] ;
   wire \r91/B[1] ;
   wire \r91/B[2] ;
   wire \r91/B[3] ;
   wire \r91/B[4] ;
   wire \r91/B[5] ;
   wire \r91/B[9] ;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire [2:0] current_state;
   wire [2:0] next_state;

   // Module instantiations
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n16),
	.SE(test_se),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.QN(n30),
	.Q(test_so),
	.D(next_state[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(deser_en),
	.B(n17),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n15),
	.A(\r91/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U8 (
	.Y(par_chk_en),
	.C(n35),
	.B(n16),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U9 (
	.Y(stp_chk_en),
	.B(n15),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n17),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U11 (
	.Y(n2),
	.B(prescale[0]),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U12 (
	.Y(next_state[2]),
	.C1(n14),
	.C0(par_error),
	.B1(n34),
	.B0(n17),
	.A1(n33),
	.A0(\r91/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n14),
	.A(par_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U14 (
	.Y(next_state[1]),
	.B1(n35),
	.B0(n36),
	.A1N(str_chk_en),
	.A0(str_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U15 (
	.Y(n36),
	.B1(n15),
	.B0(current_state[0]),
	.A1(n16),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U16 (
	.Y(str_chk_en),
	.C(n15),
	.B(current_state[1]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(next_state[0]),
	.B0(n39),
	.A1(n38),
	.A0(\r91/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U18 (
	.Y(n39),
	.B0(n41),
	.A2(par_en),
	.A1(n37),
	.A0(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U19 (
	.Y(n41),
	.D(n42),
	.C(current_state[0]),
	.B(current_state[1]),
	.A(rx_in), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U20 (
	.Y(n42),
	.B0(n30),
	.A1N(n15),
	.A0N(stp_error), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U21 (
	.Y(data_valid),
	.C(par_error),
	.B(stp_error),
	.AN(stp_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(n35),
	.B(n30),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(n40),
	.B(current_state[0]),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U24 (
	.Y(n38),
	.B(n30),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X2M U25 (
	.Y(n33),
	.C(n30),
	.B(current_state[0]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BBX1M U26 (
	.Y(n37),
	.D(bit_count[1]),
	.C(bit_count[2]),
	.BN(bit_count[0]),
	.AN(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n16),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U28 (
	.Y(n34),
	.B(n37),
	.AN(par_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U30 (
	.Y(counter_en),
	.C(n38),
	.B(n35),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U31 (
	.Y(\r91/B[0] ),
	.A(prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U32 (
	.Y(\r91/B[1] ),
	.B0(n2),
	.A1N(prescale[1]),
	.A0N(prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U33 (
	.Y(n3),
	.B(prescale[2]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U34 (
	.Y(\r91/B[2] ),
	.B0(n3),
	.A1N(prescale[2]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U35 (
	.Y(n4),
	.B(prescale[3]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U36 (
	.Y(\r91/B[3] ),
	.B0(n4),
	.A1N(prescale[3]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U37 (
	.Y(n5),
	.B(prescale[4]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U38 (
	.Y(\r91/B[4] ),
	.B0(n5),
	.A1N(prescale[4]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U39 (
	.Y(\r91/B[9] ),
	.B(prescale[5]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U40 (
	.Y(\r91/B[5] ),
	.B0(\r91/B[9] ),
	.A1(prescale[5]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U41 (
	.Y(n6),
	.B(\r91/B[0] ),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U42 (
	.Y(n9),
	.B1(n6),
	.B0(edge_count[1]),
	.A1N(\r91/B[1] ),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U43 (
	.Y(n7),
	.B(edge_count[0]),
	.AN(\r91/B[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U44 (
	.Y(n8),
	.B1(n7),
	.B0(\r91/B[1] ),
	.A1N(edge_count[1]),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BBX1M U45 (
	.Y(n13),
	.D(n8),
	.C(n9),
	.BN(\r91/B[5] ),
	.AN(\r91/B[9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n12),
	.B(edge_count[4]),
	.A(\r91/B[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n11),
	.B(edge_count[2]),
	.A(\r91/B[2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n10),
	.B(edge_count[3]),
	.A(\r91/B[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U49 (
	.Y(\r91/EQ ),
	.D(n10),
	.C(n11),
	.B(n12),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module counter_test_1 (
	clk, 
	rst, 
	counter_en, 
	prescale, 
	par_en, 
	bit_count, 
	edge_count, 
	test_si, 
	test_se, 
	FE_OFN3_SYNC_UART_SCAN_RST, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input counter_en;
   input [5:0] prescale;
   input par_en;
   output [3:0] bit_count;
   output [4:0] edge_count;
   input test_si;
   input test_se;
   input FE_OFN3_SYNC_UART_SCAN_RST;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N5;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N14;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire \add_22/carry[4] ;
   wire \add_22/carry[3] ;
   wire \add_22/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;

   // Module instantiations
   SDFFRQX2M \bit_count_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(bit_count[0]),
	.D(n38),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[3]  (
	.SI(n50),
	.SE(test_se),
	.RN(rst),
	.Q(bit_count[3]),
	.D(n36),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[2]  (
	.SI(bit_count[1]),
	.SE(test_se),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(bit_count[2]),
	.D(n46),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[1]  (
	.SI(n48),
	.SE(test_se),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(bit_count[1]),
	.D(n37),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[4]  (
	.SI(edge_count[3]),
	.SE(test_se),
	.RN(rst),
	.Q(edge_count[4]),
	.D(n42),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[3]  (
	.SI(edge_count[2]),
	.SE(test_se),
	.RN(rst),
	.Q(edge_count[3]),
	.D(n39),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[2]  (
	.SI(edge_count[1]),
	.SE(test_se),
	.RN(rst),
	.Q(edge_count[2]),
	.D(n40),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[0]  (
	.SI(n51),
	.SE(test_se),
	.RN(rst),
	.Q(edge_count[0]),
	.D(n43),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[1]  (
	.SI(n23),
	.SE(test_se),
	.RN(rst),
	.Q(edge_count[1]),
	.D(n41),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI33X2M U6 (
	.Y(n29),
	.B2(n51),
	.B1(n48),
	.B0(n33),
	.A2(n52),
	.A1(n49),
	.A0(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(n34),
	.B(n45),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n44),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n45),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U16 (
	.Y(n31),
	.C(N14),
	.B(n35),
	.A(counter_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U17 (
	.Y(n26),
	.C(n31),
	.B(n48),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U18 (
	.Y(n30),
	.B0(n31),
	.A1(n47),
	.A0(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(n35),
	.B(N12),
	.A(counter_en), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U20 (
	.Y(n37),
	.B1(n49),
	.B0(n30),
	.A1N(n26),
	.A0N(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n47),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U22 (
	.Y(n27),
	.B0(n30),
	.A1(n29),
	.A0(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U23 (
	.Y(n36),
	.B0(n25),
	.A1(n51),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U24 (
	.Y(n25),
	.D(n51),
	.C(bit_count[1]),
	.B(n26),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U25 (
	.Y(n24),
	.B0(n27),
	.A1(n50),
	.A0(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U26 (
	.Y(n2),
	.B(prescale[0]),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n46),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U28 (
	.Y(n28),
	.B1(bit_count[2]),
	.B0(n27),
	.A2(bit_count[1]),
	.A1(n50),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U29 (
	.Y(n38),
	.B1(n48),
	.B0(n45),
	.A2(n29),
	.A1(bit_count[0]),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U30 (
	.Y(n1),
	.B0N(n2),
	.A1(prescale[1]),
	.A0(prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U31 (
	.Y(n41),
	.B1(n44),
	.B0(N19),
	.A1(n34),
	.A0(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U32 (
	.Y(n40),
	.B1(n44),
	.B0(N20),
	.A1(n34),
	.A0(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U33 (
	.Y(n39),
	.B1(n44),
	.B0(N21),
	.A1(n34),
	.A0(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U34 (
	.Y(n42),
	.B1(n44),
	.B0(N22),
	.A1(n34),
	.A0(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U35 (
	.Y(n43),
	.B1(n44),
	.B0(n23),
	.A1(n34),
	.A0(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n23),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U37 (
	.Y(n32),
	.C(bit_count[3]),
	.B(n50),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(n33),
	.C(n49),
	.B(n52),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n52),
	.A(par_en), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n50),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n48),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n49),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n51),
	.A(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U44 (
	.S(N19),
	.CO(\add_22/carry[2] ),
	.B(edge_count[0]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U45 (
	.S(N20),
	.CO(\add_22/carry[3] ),
	.B(\add_22/carry[2] ),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U46 (
	.S(N21),
	.CO(\add_22/carry[4] ),
	.B(\add_22/carry[3] ),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U47 (
	.Y(N5),
	.A(prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U48 (
	.Y(n3),
	.B(prescale[2]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U49 (
	.Y(N7),
	.B0(n3),
	.A1N(prescale[2]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U50 (
	.Y(n4),
	.B(prescale[3]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U51 (
	.Y(N8),
	.B0(n4),
	.A1N(prescale[3]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U52 (
	.Y(n5),
	.B(prescale[4]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U53 (
	.Y(N9),
	.B0(n5),
	.A1N(prescale[4]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U54 (
	.Y(N11),
	.B(prescale[5]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U55 (
	.Y(N10),
	.B0(N11),
	.A1(prescale[5]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(N22),
	.B(edge_count[4]),
	.A(\add_22/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U57 (
	.Y(n22),
	.B(edge_count[3]),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U58 (
	.Y(n21),
	.B(edge_count[2]),
	.A(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U59 (
	.Y(n20),
	.B(edge_count[4]),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(n15),
	.B(N5),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U61 (
	.Y(n18),
	.B1(n1),
	.B0(n15),
	.A1(n15),
	.A0(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U62 (
	.Y(n16),
	.B(n23),
	.A(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U63 (
	.Y(n17),
	.B1(edge_count[1]),
	.B0(n16),
	.A1(n1),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U64 (
	.Y(n19),
	.D(n17),
	.C(N10),
	.B(N11),
	.AN(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U65 (
	.Y(N12),
	.D(n19),
	.C(n20),
	.B(n21),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U66 (
	.Y(N14),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampling_test_1 (
	clk, 
	rst, 
	rx_in, 
	prescale, 
	edge_count, 
	data_sample_en, 
	sampled_bit, 
	test_so, 
	test_se, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input rx_in;
   input [5:0] prescale;
   input [4:0] edge_count;
   input data_sample_en;
   output sampled_bit;
   output test_so;
   input test_se;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire sample_1;
   wire sample_2;
   wire sample_3;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire \add_34/carry[4] ;
   wire \add_34/carry[3] ;
   wire \add_34/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n14;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;

   assign test_so = sample_3 ;

   // Module instantiations
   SDFFRQX2M sample_3_reg (
	.SI(sample_2),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(sample_3),
	.D(n20),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sample_2_reg (
	.SI(sample_1),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(sample_2),
	.D(n21),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sample_1_reg (
	.SI(edge_count[4]),
	.SE(test_se),
	.RN(rst),
	.Q(sample_1),
	.D(n22),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(n17),
	.B(N12),
	.AN(data_sample_en), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n39),
	.A(rx_in), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U6 (
	.Y(n22),
	.B1(n19),
	.B0(n39),
	.A1N(sample_1),
	.A0N(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n19),
	.B(data_sample_en),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U8 (
	.Y(n21),
	.B1(n18),
	.B0(n39),
	.A1N(sample_2),
	.A0N(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U11 (
	.Y(n18),
	.B(n17),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(n20),
	.B1(n39),
	.B0(n16),
	.A1N(sample_3),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U13 (
	.Y(n16),
	.C(N20),
	.B(n17),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U14 (
	.Y(n1),
	.B(prescale[1]),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U15 (
	.S(N18),
	.CO(N19),
	.B(\add_34/carry[4] ),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U16 (
	.S(N17),
	.CO(\add_34/carry[4] ),
	.B(\add_34/carry[3] ),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U17 (
	.S(N16),
	.CO(\add_34/carry[3] ),
	.B(\add_34/carry[2] ),
	.A(prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U18 (
	.S(N15),
	.CO(\add_34/carry[2] ),
	.B(prescale[1]),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U19 (
	.Y(sampled_bit),
	.B0(n15),
	.A1N(sample_2),
	.A0N(sample_1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U20 (
	.Y(n15),
	.B0(sample_3),
	.A1(sample_2),
	.A0(sample_1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U21 (
	.Y(N6),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U22 (
	.Y(N7),
	.B0(n1),
	.A1N(prescale[2]),
	.A0N(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U23 (
	.Y(n2),
	.B(prescale[3]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U24 (
	.Y(N8),
	.B0(n2),
	.A1N(prescale[3]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U25 (
	.Y(N9),
	.B(n2),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U26 (
	.Y(N11),
	.C(n2),
	.B(prescale[5]),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U27 (
	.Y(n3),
	.B0(prescale[5]),
	.A1(n2),
	.A0(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U28 (
	.Y(N10),
	.B(n3),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U29 (
	.Y(n4),
	.B(edge_count[0]),
	.AN(N6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U30 (
	.Y(n7),
	.B1(n4),
	.B0(N7),
	.A1N(edge_count[1]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U31 (
	.Y(n5),
	.B(N6),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U32 (
	.Y(n6),
	.B1(n5),
	.B0(edge_count[1]),
	.A1N(N7),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX1M U33 (
	.Y(n14),
	.C(n6),
	.B(n7),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U34 (
	.Y(n10),
	.B(edge_count[4]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U35 (
	.Y(n9),
	.B(edge_count[2]),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(n8),
	.B(edge_count[3]),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U37 (
	.Y(N12),
	.D(n8),
	.C(n9),
	.B(n10),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n30),
	.B(edge_count[2]),
	.A(prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U39 (
	.Y(n23),
	.B(edge_count[0]),
	.AN(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U40 (
	.Y(n26),
	.B1(n23),
	.B0(prescale[2]),
	.A1N(edge_count[1]),
	.A0(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U41 (
	.Y(n24),
	.B(prescale[1]),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U42 (
	.Y(n25),
	.B1(n24),
	.B0(edge_count[1]),
	.A1N(prescale[2]),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U43 (
	.Y(n29),
	.B(n25),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U44 (
	.Y(n28),
	.B(edge_count[3]),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U45 (
	.Y(n27),
	.B(edge_count[4]),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U46 (
	.Y(N13),
	.D(n27),
	.C(n28),
	.B(n29),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U48 (
	.Y(n34),
	.B1(n4),
	.B0(N15),
	.A1N(edge_count[1]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U50 (
	.Y(n33),
	.B1(n5),
	.B0(edge_count[1]),
	.A1N(N15),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX1M U51 (
	.Y(n38),
	.C(n33),
	.B(n34),
	.AN(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n37),
	.B(edge_count[4]),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n36),
	.B(edge_count[2]),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n35),
	.B(edge_count[3]),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U55 (
	.Y(N20),
	.D(n35),
	.C(n36),
	.B(n37),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_check_test_1 (
	clk, 
	rst, 
	p_data, 
	par_typ, 
	par_chk_en, 
	sampled_bit, 
	par_error, 
	test_si, 
	test_se, 
	FE_OFN3_SYNC_UART_SCAN_RST, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input [7:0] p_data;
   input par_typ;
   input par_chk_en;
   input sampled_bit;
   output par_error;
   input test_si;
   input test_se;
   input FE_OFN3_SYNC_UART_SCAN_RST;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire par_bit;
   wire N6;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n8;
   wire n1;

   // Module instantiations
   SDFFRQX2M par_bit_reg (
	.SI(test_si),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(par_bit),
	.D(N6),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M par_error_reg (
	.SI(par_bit),
	.SE(test_se),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(par_error),
	.D(n8),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U3 (
	.Y(n8),
	.B1(par_chk_en),
	.B0(n1),
	.A1N(par_chk_en),
	.A0(par_error), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U4 (
	.Y(n1),
	.B(par_bit),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(n6),
	.B(p_data[6]),
	.A(p_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U6 (
	.Y(N6),
	.C(n4),
	.B(n3),
	.A(par_typ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U7 (
	.Y(n4),
	.C(n5),
	.B(p_data[0]),
	.A(p_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U8 (
	.Y(n3),
	.C(n6),
	.B(p_data[4]),
	.A(p_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n5),
	.B(p_data[2]),
	.A(p_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module start_check_test_1 (
	clk, 
	rst, 
	str_chk_en, 
	sampled_bit, 
	str_glitch, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input str_chk_en;
   input sampled_bit;
   output str_glitch;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;

   // Module instantiations
   SDFFRQX2M str_glitch_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(str_glitch),
	.D(n2),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U2 (
	.Y(n2),
	.B1(sampled_bit),
	.B0(str_chk_en),
	.A1N(str_chk_en),
	.A0(str_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stop_check_test_1 (
	clk, 
	rst, 
	stp_chk_en, 
	sampled_bit, 
	stp_error, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input stp_chk_en;
   input sampled_bit;
   output stp_error;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;
   wire n2;

   // Module instantiations
   SDFFRQX2M stp_error_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(stp_error),
	.D(n3),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U4 (
	.Y(n3),
	.B1(n2),
	.B0(sampled_bit),
	.A1N(n2),
	.A0N(stp_error), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n2),
	.A(stp_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_test_1 (
	clk, 
	rst, 
	deser_en, 
	sampled_bit, 
	p_data, 
	test_si, 
	test_se, 
	FE_OFN3_SYNC_UART_SCAN_RST, 
	FE_OFN12_SE, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input deser_en;
   input sampled_bit;
   output [7:0] p_data;
   input test_si;
   input test_se;
   input FE_OFN3_SYNC_UART_SCAN_RST;
   input FE_OFN12_SE;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n18;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n19;
   wire n54;
   wire [3:0] counter;

   // Module instantiations
   SDFFRQX2M \p_data_reg[5]  (
	.SI(p_data[4]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(p_data[5]),
	.D(n47),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[1]  (
	.SI(n18),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(p_data[1]),
	.D(n43),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[4]  (
	.SI(p_data[3]),
	.SE(test_se),
	.RN(rst),
	.Q(p_data[4]),
	.D(n46),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[7]  (
	.SI(p_data[6]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(p_data[7]),
	.D(n49),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[3]  (
	.SI(p_data[2]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(p_data[3]),
	.D(n45),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[6]  (
	.SI(p_data[5]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(p_data[6]),
	.D(n48),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[2]  (
	.SI(p_data[1]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(p_data[2]),
	.D(n44),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.Q(counter[3]),
	.D(n52),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(n15),
	.SE(FE_OFN12_SE),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(counter[1]),
	.D(n51),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN12_SE),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(counter[0]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(n17),
	.SE(FE_OFN8_SE),
	.RN(FE_OFN3_SYNC_UART_SCAN_RST),
	.Q(counter[2]),
	.D(n50),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \p_data_reg[0]  (
	.SI(counter[3]),
	.SE(FE_OFN8_SE),
	.RN(rst),
	.QN(n18),
	.Q(p_data[0]),
	.D(n42),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(n25),
	.B(counter[1]),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(n24),
	.B(counter[0]),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n40),
	.B(n41),
	.A(deser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(n34),
	.B(n16),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U20 (
	.Y(n51),
	.B1(n17),
	.B0(n37),
	.A1N(n25),
	.A0N(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U21 (
	.Y(n38),
	.B(n41),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n14),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n54),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n16),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U25 (
	.Y(n31),
	.C(n19),
	.B(counter[3]),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U26 (
	.Y(n49),
	.B1(n34),
	.B0(n54),
	.A1N(n34),
	.A0N(p_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U27 (
	.Y(n27),
	.B(counter[3]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U28 (
	.Y(n35),
	.B0(n37),
	.A1(n40),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U29 (
	.Y(n53),
	.B1(n40),
	.B0(counter[0]),
	.A1(n38),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U30 (
	.Y(n36),
	.B(counter[2]),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U31 (
	.Y(n45),
	.B1(n29),
	.B0(n54),
	.A1N(n29),
	.A0N(p_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n29),
	.B(n27),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U33 (
	.Y(n43),
	.B1(n26),
	.B0(n54),
	.A1N(n26),
	.A0N(p_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U34 (
	.Y(n26),
	.B(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U35 (
	.Y(n44),
	.B1(n28),
	.B0(n54),
	.A1N(n28),
	.A0N(p_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U36 (
	.Y(n28),
	.B(n27),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U37 (
	.Y(n46),
	.B1(n30),
	.B0(n54),
	.A1N(n30),
	.A0N(p_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(n30),
	.C(n31),
	.B(n17),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U39 (
	.Y(n47),
	.B1(n32),
	.B0(n54),
	.A1N(n32),
	.A0N(p_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U40 (
	.Y(n32),
	.B(n25),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U41 (
	.Y(n48),
	.B1(n33),
	.B0(n54),
	.A1N(n33),
	.A0N(p_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U42 (
	.Y(n33),
	.B(n24),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U43 (
	.Y(n50),
	.B1(n23),
	.B0(n14),
	.A1N(counter[2]),
	.A0N(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U44 (
	.Y(n52),
	.B0(n34),
	.A1N(counter[3]),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U45 (
	.Y(n39),
	.B(n35),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U46 (
	.Y(n37),
	.B0(n38),
	.A1(n40),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U47 (
	.Y(n42),
	.B(n21),
	.AN(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U48 (
	.Y(n21),
	.D(n23),
	.C(deser_en),
	.B(sampled_bit),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U49 (
	.Y(n20),
	.B0(n18),
	.A2(deser_en),
	.A1(n23),
	.A0(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U50 (
	.Y(n22),
	.D(counter[3]),
	.C(counter[2]),
	.B(n25),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U51 (
	.Y(n41),
	.D(n19),
	.C(n17),
	.B(n15),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n15),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n17),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U54 (
	.Y(n19),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U55 (
	.Y(n23),
	.B(counter[0]),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_TX_test_1 (
	CLK, 
	RST, 
	P_DATA, 
	DATA_VALID, 
	PAR_EN, 
	PAR_TYP, 
	TX_OUT, 
	BUSY, 
	test_si, 
	test_se, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] P_DATA;
   input DATA_VALID;
   input PAR_EN;
   input PAR_TYP;
   output TX_OUT;
   output BUSY;
   input test_si;
   input test_se;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PT0_;
   wire FE_UNCONNECTED_0;
   wire SER_EN;
   wire SER_DATA;
   wire SER_DONE;
   wire PAR_BIT;
   wire n3;
   wire n4;
   wire n5;
   wire [1:0] MUX_SEL;

   // Module instantiations
   serializer_WIDTH8_test_1 DUT0 (
	.CLK(CLK),
	.RST(RST),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.DATA_VALID(DATA_VALID),
	.SER_EN(SER_EN),
	.SER_DATA(SER_DATA),
	.SER_DONE(SER_DONE),
	.test_si(test_si),
	.test_so(n5),
	.test_se(test_se),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   FSM_test_1 DUT1 (
	.CLK(CLK),
	.RST(RST),
	.DATA_VALID(DATA_VALID),
	.SER_DONE(SER_DONE),
	.PAR_EN(PAR_EN),
	.SER_EN(SER_EN),
	.MUX_SEL({ MUX_SEL[1],
		MUX_SEL[0] }),
	.PAR_FLAG(FE_PT0_),
	.BUSY(BUSY),
	.test_si(n5),
	.test_so(n4),
	.test_se(test_se),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_Calc_WIDTH8_test_1 DUT2 (
	.CLK(CLK),
	.RST(RST),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.DATA_VALID(DATA_VALID),
	.PAR_TYP(PAR_TYP),
	.PAR_FLAG(SER_EN),
	.PAR_BIT(PAR_BIT),
	.test_si(n4),
	.test_so(n3),
	.test_se(test_se),
	.FE_OFN8_SE(FE_OFN8_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   MUX_test_1 DUT3 (
	.CLK(CLK),
	.RST(RST),
	.MUX_SEL({ MUX_SEL[1],
		MUX_SEL[0] }),
	.SER_DATA(SER_DATA),
	.PAR_BIT(PAR_BIT),
	.TX_OUT(TX_OUT),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module serializer_WIDTH8_test_1 (
	CLK, 
	RST, 
	P_DATA, 
	DATA_VALID, 
	SER_EN, 
	SER_DATA, 
	SER_DONE, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] P_DATA;
   input DATA_VALID;
   input SER_EN;
   output SER_DATA;
   output SER_DONE;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire [3:0] counter;
   wire [7:0] REG;

   assign test_so = counter[3] ;

   // Module instantiations
   SDFFRQX2M SER_DATA_reg (
	.SI(n52),
	.SE(test_se),
	.RN(RST),
	.Q(SER_DATA),
	.D(n39),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4]  (
	.SI(n55),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(REG[4]),
	.D(n44),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(REG[0]),
	.D(n40),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \counter_reg[3]  (
	.SN(RST),
	.SI(n18),
	.SE(FE_OFN8_SE),
	.Q(counter[3]),
	.D(n50),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \REG_reg[6]  (
	.SI(n54),
	.SE(test_se),
	.RN(RST),
	.QN(n20),
	.Q(n53),
	.D(n46),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \REG_reg[2]  (
	.SI(n57),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.QN(n23),
	.Q(n56),
	.D(n42),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \REG_reg[5]  (
	.SI(REG[4]),
	.SE(test_se),
	.RN(RST),
	.QN(n21),
	.Q(n54),
	.D(n45),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \REG_reg[1]  (
	.SI(REG[0]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.QN(n24),
	.Q(n57),
	.D(n41),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \REG_reg[7]  (
	.SI(n53),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.QN(n19),
	.Q(n52),
	.D(n47),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \REG_reg[3]  (
	.SI(n56),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.QN(n22),
	.Q(n55),
	.D(n43),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(n17),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(counter[2]),
	.D(n48),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(n16),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(counter[1]),
	.D(n49),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(SER_DATA),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(counter[0]),
	.D(n51),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n14),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U17 (
	.Y(n34),
	.B(n26),
	.A(DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n38),
	.B(n34),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U19 (
	.Y(n35),
	.B0(n36),
	.A1(n26),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U20 (
	.Y(n26),
	.B(SER_EN),
	.AN(SER_DONE), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U21 (
	.Y(n49),
	.B1(n26),
	.B0(n29),
	.A1(n17),
	.A0(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(n29),
	.B(n17),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U23 (
	.Y(n36),
	.B0(n38),
	.A1(n26),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U24 (
	.Y(n48),
	.B1(n18),
	.B0(n15),
	.A2(n29),
	.A1(counter[2]),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n15),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U26 (
	.Y(SER_DONE),
	.C(n29),
	.B(counter[3]),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U27 (
	.Y(n51),
	.B1(n26),
	.B0(counter[0]),
	.A1(n38),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U28 (
	.Y(n50),
	.B0(n34),
	.A1N(counter[3]),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(n37),
	.B(n35),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U30 (
	.Y(n41),
	.B1(n24),
	.B0(n14),
	.A1N(n14),
	.A0N(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U31 (
	.Y(n42),
	.B1(n23),
	.B0(n14),
	.A1N(n14),
	.A0N(P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U32 (
	.Y(n43),
	.B1(n22),
	.B0(n14),
	.A1N(n14),
	.A0N(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U33 (
	.Y(n45),
	.B1(n21),
	.B0(n14),
	.A1N(n14),
	.A0N(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U34 (
	.Y(n46),
	.B1(n20),
	.B0(n14),
	.A1N(n14),
	.A0N(P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U35 (
	.Y(n47),
	.B1(n19),
	.B0(n14),
	.A1N(n14),
	.A0N(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n16),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n17),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U38 (
	.Y(n40),
	.B1(n14),
	.B0(P_DATA[0]),
	.A1(REG[0]),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U39 (
	.Y(n44),
	.B1(n14),
	.B0(P_DATA[4]),
	.A1(REG[4]),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U40 (
	.Y(n30),
	.B1(n31),
	.B0(counter[1]),
	.A2(REG[4]),
	.A1(n17),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U41 (
	.Y(n31),
	.B1(n21),
	.B0(counter[0]),
	.A1(n20),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U42 (
	.Y(n32),
	.B1(n33),
	.B0(counter[1]),
	.A2(counter[0]),
	.A1(n17),
	.A0(REG[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U43 (
	.Y(n33),
	.B1(n24),
	.B0(counter[0]),
	.A1(n23),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U44 (
	.Y(n39),
	.B1(n26),
	.B0(n25),
	.A1N(n26),
	.A0N(SER_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U45 (
	.Y(n25),
	.B1(n28),
	.B0(counter[2]),
	.A1(n18),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U46 (
	.Y(n27),
	.B0(n32),
	.A1(n19),
	.A0(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U47 (
	.Y(n28),
	.B0(n30),
	.A1(n22),
	.A0(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n18),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_test_1 (
	CLK, 
	RST, 
	DATA_VALID, 
	SER_DONE, 
	PAR_EN, 
	SER_EN, 
	MUX_SEL, 
	PAR_FLAG, 
	BUSY, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input DATA_VALID;
   input SER_DONE;
   input PAR_EN;
   output SER_EN;
   output [1:0] MUX_SEL;
   output PAR_FLAG;
   output BUSY;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n5;
   wire n6;
   wire n11;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n5),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n11),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U6 (
	.Y(BUSY),
	.B(n10),
	.AN(SER_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(next_state[2]),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U8 (
	.Y(next_state[0]),
	.C(current_state[0]),
	.B(current_state[2]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U9 (
	.Y(n9),
	.B1(n11),
	.B0(DATA_VALID),
	.A2(PAR_EN),
	.A1(current_state[1]),
	.A0(SER_DONE), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U10 (
	.Y(n8),
	.B(current_state[1]),
	.AN(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n5),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U12 (
	.Y(next_state[1]),
	.B1(n6),
	.B0(n8),
	.A2(current_state[1]),
	.A1(current_state[2]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U14 (
	.Y(n7),
	.B0(current_state[0]),
	.A1N(PAR_EN),
	.A0(SER_DONE), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U15 (
	.Y(n10),
	.C(current_state[2]),
	.B(n11),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n11),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(MUX_SEL[0]),
	.B0(n10),
	.A1(n8),
	.A0(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U18 (
	.Y(MUX_SEL[1]),
	.B0(n10),
	.A1(n5),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U20 (
	.Y(SER_EN),
	.B0(n8),
	.A1(n5),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_Calc_WIDTH8_test_1 (
	CLK, 
	RST, 
	P_DATA, 
	DATA_VALID, 
	PAR_TYP, 
	PAR_FLAG, 
	PAR_BIT, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN8_SE, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] P_DATA;
   input DATA_VALID;
   input PAR_TYP;
   input PAR_FLAG;
   output PAR_BIT;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN8_SE;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n10;
   wire n11;
   wire n12;
   wire [7:0] REG;

   assign test_so = REG[7] ;

   // Module instantiations
   SDFFRQX2M PAR_BIT_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(PAR_BIT),
	.D(n21),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[5]  (
	.SI(REG[4]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[5]),
	.D(n27),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[1]  (
	.SI(REG[0]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(REG[1]),
	.D(n23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[4]  (
	.SI(REG[3]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[4]),
	.D(n26),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[0]  (
	.SI(PAR_BIT),
	.SE(test_se),
	.RN(RST),
	.Q(REG[0]),
	.D(n22),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[2]  (
	.SI(REG[1]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(REG[2]),
	.D(n24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[3]  (
	.SI(REG[2]),
	.SE(FE_OFN8_SE),
	.RN(RST),
	.Q(REG[3]),
	.D(n25),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[6]  (
	.SI(REG[5]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[6]),
	.D(n28),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \REG_reg[7]  (
	.SI(REG[6]),
	.SE(test_se),
	.RN(RST),
	.Q(REG[7]),
	.D(n29),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n12),
	.A(PAR_FLAG), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U13 (
	.Y(n20),
	.B(n12),
	.A(DATA_VALID), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n11),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n14),
	.B(n12),
	.A(PAR_TYP), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U16 (
	.Y(n21),
	.B0(n13),
	.A1N(n12),
	.A0N(PAR_BIT), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U17 (
	.Y(n13),
	.B1(n15),
	.B0(n14),
	.A2(n10),
	.A1(n11),
	.A0(PAR_FLAG), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n10),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U19 (
	.Y(n15),
	.B(n17),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U20 (
	.Y(n22),
	.B1(n20),
	.B0(P_DATA[0]),
	.A1N(n20),
	.A0(REG[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U21 (
	.Y(n23),
	.B1(n20),
	.B0(P_DATA[1]),
	.A1N(n20),
	.A0(REG[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U22 (
	.Y(n24),
	.B1(n20),
	.B0(P_DATA[2]),
	.A1N(n20),
	.A0(REG[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U23 (
	.Y(n25),
	.B1(n20),
	.B0(P_DATA[3]),
	.A1N(n20),
	.A0(REG[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U24 (
	.Y(n26),
	.B1(n20),
	.B0(P_DATA[4]),
	.A1N(n20),
	.A0(REG[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U25 (
	.Y(n27),
	.B1(n20),
	.B0(P_DATA[5]),
	.A1N(n20),
	.A0(REG[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U26 (
	.Y(n28),
	.B1(n20),
	.B0(P_DATA[6]),
	.A1N(n20),
	.A0(REG[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U27 (
	.Y(n29),
	.B1(n20),
	.B0(P_DATA[7]),
	.A1N(n20),
	.A0(REG[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U28 (
	.Y(n17),
	.C(n18),
	.B(REG[4]),
	.A(REG[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U29 (
	.Y(n18),
	.B(REG[6]),
	.A(REG[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U30 (
	.Y(n16),
	.C(n19),
	.B(REG[0]),
	.A(REG[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U31 (
	.Y(n19),
	.B(REG[3]),
	.A(REG[2]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module MUX_test_1 (
	CLK, 
	RST, 
	MUX_SEL, 
	SER_DATA, 
	PAR_BIT, 
	TX_OUT, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [1:0] MUX_SEL;
   input SER_DATA;
   input PAR_BIT;
   output TX_OUT;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N13;
   wire n2;

   // Module instantiations
   SDFFSQX2M TX_OUT_reg (
	.SN(RST),
	.SI(test_si),
	.SE(test_se),
	.Q(TX_OUT),
	.D(N13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U5 (
	.Y(N13),
	.B0(n2),
	.A1N(MUX_SEL[0]),
	.A0N(SER_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U6 (
	.Y(n2),
	.B0(MUX_SEL[1]),
	.A1(PAR_BIT),
	.A0(MUX_SEL[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_TOP (
	scan_clk, 
	scan_rst, 
	test_mode, 
	SE, 
	SI, 
	SO, 
	REF_CLK, 
	RST, 
	UART_CLK, 
	RX_IN, 
	TX_OUT, 
	PARITY_ERROR, 
	STOP_ERROR, 
	BUSY, 
	VDD, 
	VSS);
   input scan_clk;
   input scan_rst;
   input test_mode;
   input SE;
   input [3:0] SI;
   output [3:0] SO;
   input REF_CLK;
   input RST;
   input UART_CLK;
   input RX_IN;
   output TX_OUT;
   output PARITY_ERROR;
   output STOP_ERROR;
   output BUSY;
   inout VDD;
   inout VSS;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L7_N0;
   wire scan_clk__L6_N1;
   wire scan_clk__L6_N0;
   wire scan_clk__L5_N1;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N1;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire REF_SCAN_CLK__L2_N1;
   wire REF_SCAN_CLK__L2_N0;
   wire REF_SCAN_CLK__L1_N0;
   wire UART_SCAN_CLK__L6_N0;
   wire UART_SCAN_CLK__L5_N0;
   wire UART_SCAN_CLK__L4_N1;
   wire UART_SCAN_CLK__L4_N0;
   wire UART_SCAN_CLK__L3_N1;
   wire UART_SCAN_CLK__L3_N0;
   wire UART_SCAN_CLK__L2_N1;
   wire UART_SCAN_CLK__L2_N0;
   wire UART_SCAN_CLK__L1_N1;
   wire UART_SCAN_CLK__L1_N0;
   wire UART_RX_SCAN_CLK__L1_N0;
   wire UART_TX_SCAN_CLK__L1_N0;
   wire FE_OFN12_SE;
   wire FE_OFN10_SE;
   wire FE_OFN9_SE;
   wire FE_OFN8_SE;
   wire FE_OFN7_SE;
   wire FE_OFN6_SE;
   wire FE_OFN3_SYNC_UART_SCAN_RST;
   wire FE_OFN1_SYNC_REF_SCAN_RST;
   wire FE_OFN0_SYNC_REF_SCAN_RST;
   wire REF_SCAN_CLK;
   wire UART_SCAN_CLK;
   wire RX_CLK;
   wire UART_RX_SCAN_CLK;
   wire TX_CLK;
   wire UART_TX_SCAN_CLK;
   wire RSTN_SCAN_RST;
   wire REF_SYNC_RST;
   wire SYNC_REF_SCAN_RST;
   wire UART_SYNC_RST;
   wire SYNC_UART_SCAN_RST;
   wire RX_DATA_VALID;
   wire SYNC_RX_DATA_VALID;
   wire RD_DATA_VALID;
   wire ALU_OUT_VALID;
   wire FIFO_FULL;
   wire ALU_EN;
   wire CLK_GATE_EN;
   wire WR_EN;
   wire RD_EN;
   wire CTRL_OUT_VALID;
   wire _0_net_;
   wire ALU_CLK;
   wire RD_INC;
   wire FIFO_EMPTY;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n11;
   wire n12;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n22;
   wire n23;
   wire n24;
   wire [7:0] RX_P_DATA;
   wire [7:0] SYNC_RX_P_DATA;
   wire [7:0] RD_DATA;
   wire [15:0] ALU_OUT;
   wire [3:0] FUN;
   wire [3:0] ADDRESS;
   wire [7:0] WR_DATA;
   wire [7:0] CTRL_OUT_DATA;
   wire [7:0] OP_A;
   wire [7:0] OP_B;
   wire [7:0] UART_config;
   wire [7:0] TX_DIV_RATIO;
   wire [7:0] RX_DIV_RATIO;
   wire [7:0] TX_IN_DATA;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;
   wire SYNOPSYS_UNCONNECTED__3;

   assign SO[2] = UART_config[2] ;
endmodule

